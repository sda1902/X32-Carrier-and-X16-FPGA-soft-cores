module EU64X16E (
	input wire CLK, RESET, CLOAD,
	input wire [7:0] CPU,
	input wire [15:0] TASKID,
	input wire [23:0] CPSR,
	// interface to datapatch of memory subsystem
	input wire NEXT, StreamNEXT, NetNEXT,
	output reg ACT, StreamACT, NetACT, CMD, 
	output reg [1:0] OS,
	output reg [44:0] ADDRESS,
	output reg [36:0] OFFSET,
	output reg [31:0] SELECTOR,
	output reg [63:0] DTo,
	output reg [7:0] TAGo,
	input wire DRDY,
	input wire [7:0] TAGi,
	input wire [2:0] SZi,
	input wire [63:0] DTi,
	// FFT memory interface
	input wire FFTMemNEXT, FFTNetNEXT,
	output wire FFTMemACT, FFTNetACT, FFTMemCMD,
	output wire [41:0] FFTMemADDR,
	output wire [33:0] FFTMemOFFSET,
	output wire [31:0] FFTMemSEL,
	output wire [63:0] FFTMemDO,
	output wire [7:0] FFTMemTO,
	// interface to the descriptor pre-loading system
	input wire [39:0] DTBASE,
	input wire [23:0] DTLIMIT,
	input wire [1:0] CPL,
	// interface to message control subsystem
	output wire [63:0] PARAM,
	output wire [3:0] PARREG,
	output wire MSGREQ, MALLOCREQ, PARREQ, ENDMSG, BKPT,
	output reg EMPTY,
	output wire HALT,
	output wire NPCS,
	output wire SMSGBKPT,
	input wire CEXEC, ESMSG, CONTINUE,
	input wire CSTOP, LIRESET,
	// context store interface
	input wire [5:0] RA,
	output reg [63:0] CDATA,
	output wire [36:0] RIP,
	// error reporting interface
	output wire ESTB,
	output wire [28:0] ECD,
	// FFT engine error report interface
	output wire FFTESTB,
	output wire [28:0] FFTECD,
	output wire [23:0] FFTCPSR,
	// test purpose pins
	output wire FATAL,
	// Performance monitor outputs
	output reg [3:0] IV,
	output wire [23:0] CSEL
	);

integer i;

// general purpose register file
reg [127:0] GPR [15:0];
// arithmetic flags
reg [31:0] AFR [15:0];
reg [15:0] FlagWrite;
reg ContextLoadFlag;
// address register file
reg [36:0] ADR [15:0];
// GPR valid flags
reg [15:0] GPVFReg;
wire [15:0] GPVFINVD;

// FACC unit resources
wire [19:0] FMULACCBus;
reg [19:0] FMULACCReg; //0 - ACT, 3:1 - ctrlSel, 7:4 - DST, 11:8 - CtrlOffsetReg, 15:12 - DataOffsetReg, 18:16 - DataSel, 19-CMD
reg FMULACCACTReg, FMULACCCMDReg, FFT32NEXTReg;
wire FMULACCNEXT;
reg [3:0] FMULACCDSTReg;
reg [2:0] FMULACCDataSelReg, FMULACCCtrlSelReg;
reg [34:0] FMULACCDataOffsetReg;
reg [33:0] FMULACCCtrlOffsetReg;
wire FMULACCRDY, FMULACCSIGN, FMULACCZERO, FMULACCINF, FMULACCNAN;
wire [31:0] FMULACCR;
wire [3:0] FMULACCDST;
wire FMULACCMemACT, FMULACCSIZE, FMULACCTAGo;
wire [2:0] FMULACCMemSEL;
wire [34:0] FMULACCMemOffset;
reg FMULACCDRDYFlag;
reg [9:0] FMULACCBypassControlOffsetReg, FMULACCBypassDataOffsetReg, FFTBypassReg;
wire SkipFifoData, SkipFifoFlag;
reg [4:0] FFTParReg;

// FFT resources
wire FFT32NEXT;
reg [31:0] FFTDataSelReg, FFTCtrlSelReg;
reg [33:0] FFTDataBaseReg, FFTCtrlBaseReg;
reg [18:0] FFTIndexReg;

// FADD unit resources
wire [13:0] FADDInstBusA, FADDInstBusB;
reg [13:0] FADDInstRegA, FADDInstRegB;
reg [127:0] FADDARegA, FADDBRegA, FADDARegB, FADDBRegB;
reg [2:0] FADDSARegA, FADDSBRegA, FADDSARegB, FADDSBRegB;
reg [3:0] FADDDSTRegA, FADDDSTRegB, FADDDSTRA, FADDDSTRB;
reg [9:0] FADDBypassARegA, FADDBypassARegB, FADDBypassBRegA, FADDBypassBRegB;
reg FADDACTRegA, FADDCMDRegA, FADDACTRegB, FADDCMDRegB, FADDRDYRA, FADDRDYRB;
wire [127:0] FADDRA, FADDRB;
wire [3:0] FADDDSTA, FADDDSTB;
wire [2:0] FADDSRA, FADDSRB;
wire FADDRDYA, FADDZeroA, FADDSignA, FADDInfA, FADDNaNA, FADDRDYB, FADDZeroB, FADDSignB, FADDInfB, FADDNaNB;

// FMUL resources
wire [12:0] FMULInstBusA, FMULInstBusB;
reg [12:0] FMULInstRegA, FMULInstRegB;
reg [127:0] FMULARegA, FMULBRegA, FMULARegB, FMULBRegB;
reg FMULACTRegA, FMULACTRegB;
reg [2:0] FMULSARegA, FMULSBRegA, FMULSARegB, FMULSBRegB;
reg [3:0] FMULDSTRegA, FMULDSTRegB;
reg [9:0] FMULBypassARegA, FMULBypassARegB, FMULBypassBRegA, FMULBypassBRegB;
wire [63:0] FMULRA, FMULRB;
wire [127:0] FMULRQA, FMULRQB;
wire [3:0] FMULDSTA [1:0];
wire [3:0] FMULDSTB [1:0];
wire FMULSRA, FMULSRB;
wire [1:0] FMULRDYA, FMULZeroA, FMULSignA, FMULInfA, FMULNaNA, FMULRDYB, FMULZeroB, FMULSignB, FMULInfB, FMULNaNB;
reg [1:0] FMULRDYRA, FMULRDYRB;
reg [3:0] FMULDSTRA [1:0];
reg [3:0] FMULDSTRB [1:0];

// FDIV unit resources
wire [13:0] FDIVInstBus;
reg [13:0] FDIVInstReg;
reg [127:0] FDIVAReg, FDIVBReg;
reg FDIVACTReg, FDIVCMDReg;
reg [2:0] FDIVSAReg, FDIVSBReg, FDIVSRReg;
reg [3:0] FDIVDSTReg;
reg [9:0] FDIVBypassAReg, FDIVBypassBReg;
wire [127:0] FDIVR;
wire [3:0] FDIVDST;
wire [2:0] FDIVSR;
wire FDIVRDY, FDIVZero, FDIVInf, FDIVNaN, FDIVSign, FDIVNEXT;

// Integer ALU Resources
wire [24:0] ALUInstBusA, ALUInstBusB;
reg [24:0] ALUInstRegA, ALUInstRegB;
reg ALUACTRegA, ALUACTRegB, ALURDYRA, ALURDYRB;
reg [63:0] ALUARegA, ALUBRegA, ALUCRegA, ALUDRegA, ALUARegB, ALUBRegB, ALUCRegB, ALUDRegB;
reg [1:0] ALUSARegA, ALUSBRegA, ALUSCRegA, ALUSDRegA, ALUSRRegA, ALUSARegB, ALUSBRegB, ALUSCRegB, ALUSDRegB, ALUSRRegB;
reg [2:0] ALUOpCODERegA, ALUOpCODERegB;
reg [3:0] ALUDSTRegA, ALUDSTRegB, ALUDSTRA, ALUDSTRB;
reg [9:0] ALUBypassARegA, ALUBypassBRegA, ALUBypassCRegA, ALUBypassDRegA, ALUBypassARegB, ALUBypassBRegB, ALUBypassCRegB, ALUBypassDRegB;
wire [63:0] ALURA, ALURB;
wire [3:0] ALUDSTA, ALUDSTB;
wire ALURDYA, ALUOVRA, ALUSignA, ALUZeroA, ALURDYB, ALUOVRB, ALUSignB, ALUZeroB;
wire [15:0] ALUCOUTA, ALUCOUTB;
wire [1:0] ALUSRA, ALUSRB;

// Parallel shifter resources
wire [12:0] ShiftInstBus;
reg [12:0] ShiftInstReg;
reg [63:0] ShiftAReg;
reg [5:0] ShiftBReg;
reg [9:0] ShiftBypassAReg, ShiftBypassBReg;
reg [3:0] ShiftDSTReg, ShiftDSTR;
reg [2:0] ShiftOPRReg;
reg [1:0] ShiftSAReg, ShiftSRReg;
reg ShiftACTReg, ShiftRDYR;
wire [63:0] ShiftR;
wire [3:0] ShiftDST;
wire ShiftRDY, ShiftOVR, ShiftZERO, ShiftCOUT, ShiftSign;
wire [1:0] ShiftSR;

// miscellaneous unit resources
wire [11:0] MiscInstBus;
reg [11:0] MiscInstReg;
reg [2:0] MiscOPRReg;
reg MiscACTReg, MiscRDYR;
reg [127:0] MiscAReg;
reg [3:0] MiscDSTReg, MiscDSTR;
reg [2:0] MiscSAReg, MiscSDReg, MiscSRReg;
reg [15:0] MiscCINReg;
reg [9:0] MiscBypassAReg, MiscBypassBReg;
wire [127:0] MiscR;
wire [3:0] MiscDST;
wire [2:0] MiscSR;
wire MiscRDY, MiscCOUT, MiscOVR, MiscSign, MiscZero, MiscNaN;

// data movement resources
reg [14:0] MovInstReg;
wire [14:0] MovInstBus;
reg [127:0] MovReg;
reg [2:0] MovSR;
reg [15:0] LIResetFlag, LIFlag;
reg [9:0] CopyBypassReg;

// loop instruction bus
reg [15:0] LoopInstReg;
wire [15:0] LoopInstBus;
reg LoopInstFlag;
reg [9:0] LoopBypassReg;

// prefetch control resources
reg [16:0] PrefInstReg;
wire [16:0] PrefInstBus;
reg [9:0] PrefBypassReg, PrefCCBypassReg;
wire IFetch, InsRDY, PrefACT, PrefCall, PrefRet, PrefEMPTY, PrefERST, CodeError;
wire [3:0] IVF;
wire [63:0] INST;
wire [36:0] PrefOffset;
wire [35:0] PrefRealIP;
wire [2:0] PrefTag;
reg PrefCC, PrefCallReg, PrefRetReg;
wire SeqEMPTY, MFLag;

// memory read/write resources
reg [15:0] MemInstReg;
wire [15:0] MemInstBus;
reg MemDelayFlag, MemFifoFullFlag;
wire [216:0] MemFifoBus;
wire MemFifoEmpty;
wire [5:0] MemFifoUsedW;
reg MemBusy, MemReq, MemLoadSel, MemOpr, MemADRPushPop, MemPUSH, MemPOP, MemLDST, MemLDO, MemLoadOffset, MemSecondCycle, MemReadAR, MemLSelNode, MemNext;
reg [2:0] MemSEL, MemSize, MemAMode;
reg [31:0] MemAFR;
reg [36:0] ARData, MemGPROffset;
reg [127:0] MemGPR;
reg [3:0] MemDST, MemOFF;
reg [4:0] MemoryOSValue;
reg [15:0] MemASelNode, MemFSelNode;
reg [1:0] MemCNT;
reg [2:0] SZiReg;
reg [7:0] TAGiReg;

// check memory access stage
reg CheckACT, CheckCMD, CheckNetwork, CheckNext, CheckPref;
reg [1:0] CheckOS;
reg [36:0] CheckOffset;
reg [31:0] CheckLL, CheckUL, CheckSelector;
reg [3:0] CheckAR;
reg [39:0] CheckBase;
reg [23:0] CheckLowerSel, CheckUpperSel;
reg [63:0] CheckData;
reg [7:0] CheckTag;
reg [2:0] CheckSEL;

/*
descriptor registers
39:0	- base address		40
71:40	- lower limit		32
103:72	- upper limit		32
127:104	- lower selector	24
151:128 - upper selector	24
154:152 - access rights		4
155 	- valid bit
*/
reg [155:0] DTR [7:0];
reg [8:0] DTRWriteFlag;
reg DTRLoadedFlag, DescriptorLoadState, ValidDescriptor, LoadNewDSC, LoadLowerDSC, LoadUpperDSC, RetryTransactionFlag;
reg [23:0] DLSelector;
// state machine for descriptor loading
reg [3:0] DLMachine;
parameter WS=4'd0, CSS=4'd1, ZSS=4'd2, INVSS=4'd3, LBS=4'd4, LLSS=4'd5, LSLS=4'd6, RWS=4'd7, INVOBS=4'd8, STS=4'd9, AERSS=4'd10;
reg SkipDataRead, InvalidType, InvalidCPL, InvalidTaskID, AccessError;
reg [3:0] STAGReg;
reg [23:0] InvalidSelector;


// wire result flags
reg [15:0] GPRByteNode, GPRWordNode, GPRDwordNode, GPRQwordNode, GPROwordNode, FADDSelNodeA, FADDSelNodeB, FMULSelNodeA, FMULQSelNodeA, FMULSelNodeB, FMULQSelNodeB, 
			FMULACCSelNode, FDIVSelNode, ALUSelNodeA, ALUSelNodeB, ShiftSelNode, MiscSelNode, MovSelNode, MemSelNode, MemARSelNode,
			FFTSelNode;

/*
===========================================================================================================
				Modules
===========================================================================================================
*/
// memory operations queue														55							54:52						51:15				14:0
sc_fifo MemFIFO (.data({PrefRet, PrefCall, AFR[MemInstReg[15:12]], PrefCall ? {91'd0,PrefRealIP,1'b0}:GPR[MemInstReg[15:12]], AFR[MemInstReg[11:8]][27:25], GPR[MemInstReg[11:8]][36:0], MemInstReg[15:1]}),
				.wrreq((MemInstReg[0] & ~MemDelayFlag & ~MemFifoFullFlag) | PrefCall | PrefRet),
				.rdreq((~MemBusy | (MemNext & ~FMULACCMemACT) | MemLoadOffset | (MemLoadSel & (MemDST!={CheckSEL,CheckACT})) | MemReadAR) & ~MemCNT[1] & ~MemCNT[0]),
				.clock(CLK), .sclr(~RESET), .q(MemFifoBus), .empty(MemFifoEmpty), .almost_empty(), .usedw(MemFifoUsedW));
defparam MemFIFO.LPM_WIDTH=217, MemFIFO.LPM_NUMWORDS=64, MemFIFO.LPM_WIDTHU=6;
 
// Instruction prefetcher
PrefetcherX16 Pref (.CLK(CLK), .RESET(RESET), .CSELCHG(MemASelNode[13]), .DRDY(DRDY), .TAGi(TAGi), .DTi(DTi), .IFETCH(IFetch), .IRDY(InsRDY),
				.VF(IVF), .IBUS(INST), .NEXT(~MemReq & MemNext & ~FMULACCMemACT & ~PrefCallReg & ~PrefRetReg), .ACT(PrefACT), .OFFSET(PrefOffset), .TAGo(PrefTag),
				// instruction for prefetcher
				.CBUS(LoopInstFlag ? {LoopInstReg, 1'b1} : PrefInstReg),
				.GPRBUS(LoopInstFlag ? ((GPR[LoopInstReg[15:12]][63:0] & {64{~(|LoopBypassReg)}}) |
										(FADDRA[63:0] & {64{LoopBypassReg[0]}}) |
										(FMULRA & {64{LoopBypassReg[1]}}) |
										(FMULRQA[63:0] & {64{LoopBypassReg[2]}}) |
										(ALURA & {64{LoopBypassReg[3]}}) |
										(ShiftR & {64{LoopBypassReg[4]}}) |
										(MiscR[63:0] & {64{LoopBypassReg[5]}}) |
										(FADDRB[63:0] & {64{LoopBypassReg[6]}}) |
										(FMULRB & {64{LoopBypassReg[7]}}) |
										(FMULRQB[63:0] & {64{LoopBypassReg[8]}}) |
										(ALURB & {64{LoopBypassReg[9]}})) :
									   ((GPR[PrefInstReg[16:13]][63:0] & {64{~(|PrefBypassReg)}}) |
										(FADDRA[63:0] & {64{PrefBypassReg[0]}}) |
										(FMULRA & {64{PrefBypassReg[1]}}) |
										(FMULRQA[63:0] & {64{PrefBypassReg[2]}}) |
										(ALURA & {64{PrefBypassReg[3]}}) |
										(ShiftR & {64{PrefBypassReg[4]}}) |
										(MiscR[63:0] & {64{PrefBypassReg[5]}}) |
										(FADDRB[63:0] & {64{PrefBypassReg[6]}}) |
										(FMULRB & {64{PrefBypassReg[7]}}) |
										(FMULRQB[63:0] & {64{PrefBypassReg[8]}}) |
										(ALURB & {64{PrefBypassReg[9]}}))),
				// flags
				.CC(PrefCC), .MOVFLAG(MFLag | MemInstReg[0]), .CALL(PrefCall), .RET(PrefRet), .ERST(PrefERST), .RIP(PrefRealIP), .CEXEC(CEXEC),
				.ESMSG(ESMSG), .CONTINUE(CONTINUE), .STOP(CSTOP | ESTB),
				// interface to message and memory control system
				.GPINDX(PARREG),
				.SMSG(MSGREQ), .MALLOC(MALLOCREQ), .GPAR(PARREQ), .EMSG(ENDMSG), .BKPT(BKPT), .EMPTY(PrefEMPTY), .HALT(HALT), .PARAM(PARAM),
				.SLEEP(NPCS), .SMSGBKPT(SMSGBKPT),
				// code fetch error
				.CFERROR(CodeError),
				// Fatal error reporting
				.FATAL(FATAL)
				);


// Instruction sequencer
SequencerX16E Seq (.CLK(CLK), .RESET(RESET), .IRDY(InsRDY), .VF(IVF), .IBUS(INST),
				.IRD(IFetch), .GPRVF(GPVFReg), .GPRINVD(GPVFINVD), .EMPTY(SeqEMPTY), .MOVFLAG(MFLag), .FDIVRDY(~FDIVInstReg[0]), .FMULACCRDY(~FMULACCReg[0]),
				.MEMRDY(~MemDelayFlag & ~MemFifoFullFlag), .FADDBusA(FADDInstBusA), .FADDBusB(FADDInstBusB), .FMULBusA(FMULInstBusA), .FMULBusB(FMULInstBusB),
				.FMULACCBus(FMULACCBus), .FDIVBus(FDIVInstBus), .ALUBusA(ALUInstBusA), .ALUBusB(ALUInstBusB), .ShiftBus(ShiftInstBus),
				.MiscBus(MiscInstBus), .LoopBus(LoopInstBus), .MovBus(MovInstBus), .MemBus(MemInstBus), .CtrlBus(PrefInstBus));

// 32-bit multiplier/accumulator
Neuro16 FMULACC (.CLK(CLK), .RESET(RESET), .ACT(FMULACCACTReg & ~FMULACCCMDReg), .MAERR(CheckACT & CheckCMD & (DLMachine==STS) & (CheckTag[7:1]==7'b1100000)),
				.NEXT(FMULACCNEXT), .DSTi(FMULACCDSTReg), .DataSEL(FMULACCDataSelReg), .CtrlSEL(FMULACCCtrlSelReg), .DataOffset(FMULACCDataOffsetReg),
				.CtrlOffset(FMULACCCtrlOffsetReg), .RDY(FMULACCRDY), .SIGN(FMULACCSIGN), .ZERO(FMULACCZERO), .INF(FMULACCINF), .NAN(FMULACCNAN),
				.R(FMULACCR), .DSTo(FMULACCDST),
				// memory interface
				.MemNEXT(MemNext), .MemACT(FMULACCMemACT), .MemSEL(FMULACCMemSEL), .MemOffset(FMULACCMemOffset), .SIZE(FMULACCSIZE),
				.TAGo(FMULACCTAGo), .DRDY(FMULACCDRDYFlag | SkipFifoFlag),
				.TAGi((TAGiReg[0] & FMULACCDRDYFlag) | (SkipFifoData & ~FMULACCDRDYFlag)), .DTi(DTi));

SFifo SkipFifo(.CLK(CLK), .RST(RESET), .D(CheckTag[0]), .WR(CheckACT & CheckCMD & (DLMachine==STS) & (CheckTag[7:1]==7'b1100000)),
				.Q(SkipFifoData), .VALID(SkipFifoFlag), .RD(~FMULACCDRDYFlag));


// 32-bit FFT processor
fftX16 FFT32(.CLK(CLK), .RESET(RESET), .CPU(CPU), .DTBASE(DTBASE), .DTLIMIT(DTLIMIT), .CPL(CPL), .TASKID(TASKID), .CPSR(CPSR),
				// command interface
				.NEXT(FFT32NEXT), .ACT(FMULACCACTReg & FMULACCCMDReg), .DataObject(FFTDataSelReg), .ControlObject(FFTCtrlSelReg),
				.DataOffset(FFTDataBaseReg+FMULACCDataOffsetReg[34:1]), .ControlOffset(FFTCtrlBaseReg+FMULACCCtrlOffsetReg),
				.PAR(FFTParReg), .INDEX(FFTIndexReg),
				// memory interface
				.MemNEXT(FFTMemNEXT), .NetNEXT(FFTNetNEXT), .MemACT(FFTMemACT), .NetACT(FFTNetACT), .MemCMD(FFTMemCMD), .MemADDR(FFTMemADDR),
				.MemOFFSET(FFTMemOFFSET), .MemSEL(FFTMemSEL), .MemDO(FFTMemDO), .MemTO(FFTMemTO), .MemDRDY(DRDY), .MemDI(DTi), .MemTI(TAGi),
				// error report interface
				.ESTB(FFTESTB), .ECD(FFTECD), .ECPSR(FFTCPSR));
				
// 128-bit adder modules
FPADD128 FPAdderA(.CLK(CLK), .RESET(RESET), .ACT(FADDACTRegA), .CMD(FADDCMDRegA), .A(FADDARegA), .B(FADDBRegA),
		.SA(FADDSARegA), .SB(FADDSBRegA), .DSTI(FADDDSTRegA), .RDY(FADDRDYA), .SIGN(FADDSignA), .ZERO(FADDZeroA), .INF(FADDInfA),
		.NAN(FADDNaNA), .SR(FADDSRA), .DSTO(FADDDSTA), .R(FADDRA));
FPADD128 FPAdderB(.CLK(CLK), .RESET(RESET), .ACT(FADDACTRegB), .CMD(FADDCMDRegB), .A(FADDARegB), .B(FADDBRegB),
		.SA(FADDSARegB), .SB(FADDSBRegB), .DSTI(FADDDSTRegB), .RDY(FADDRDYB), .SIGN(FADDSignB), .ZERO(FADDZeroB), .INF(FADDInfB),
		.NAN(FADDNaNB), .SR(FADDSRB), .DSTO(FADDDSTB), .R(FADDRB));

// 128-bit FP multiplier
FPMUL128 FPMultA (.CLK(CLK), .RESET(RESET), .ACT(FMULACTRegA), .DSTI(FMULDSTRegA), .A(FMULARegA), .B(FMULBRegA),
				.SA(FMULSARegA), .SB(FMULSBRegA), .RDYSD(FMULRDYA[0]), .RDYQ(FMULRDYA[1]), .ZEROSD(FMULZeroA[0]), .SIGNSD(FMULSignA[0]),
				.INFSD(FMULInfA[0]), .NANSD(FMULNaNA[0]), .ZEROQ(FMULZeroA[1]), .SIGNQ(FMULSignA[1]), .INFQ(FMULInfA[1]),
				.NANQ(FMULNaNA[1]), .SR(FMULSRA), .DSTSD(FMULDSTA[0]), .DSTQ(FMULDSTA[1]), .RSD(FMULRA), .RQ(FMULRQA));
FPMUL128 FPMultB (.CLK(CLK), .RESET(RESET), .ACT(FMULACTRegB), .DSTI(FMULDSTRegB), .A(FMULARegB), .B(FMULBRegB),
				.SA(FMULSARegB), .SB(FMULSBRegB), .RDYSD(FMULRDYB[0]), .RDYQ(FMULRDYB[1]), .ZEROSD(FMULZeroB[0]), .SIGNSD(FMULSignB[0]),
				.INFSD(FMULInfB[0]), .NANSD(FMULNaNB[0]), .ZEROQ(FMULZeroB[1]), .SIGNQ(FMULSignB[1]), .INFQ(FMULInfB[1]),
				.NANQ(FMULNaNB[1]), .SR(FMULSRB), .DSTSD(FMULDSTB[0]), .DSTQ(FMULDSTB[1]), .RSD(FMULRB), .RQ(FMULRQB));

// FP 64-bit divisor
FPDIV128 FDIV (.CLK(CLK), .ACT(FDIVACTReg), .CMD(FDIVCMDReg), .SA(FDIVSAReg), .SB(FDIVSBReg), .RST(RESET), .A(FDIVAReg), .B(FDIVBReg),
				.DSTi(FDIVDSTReg), .R(FDIVR), .DSTo(FDIVDST), .RDY(FDIVRDY), .Zero(FDIVZero), .Inf(FDIVInf),
				.NaN(FDIVNaN), .Sign(FDIVSign), .SR(FDIVSR), .NEXT(FDIVNEXT));

// integer ALU
ALU64X16 IntALUA (.CLK(CLK), .ACT(ALUACTRegA), .CIN(1'b0), .DSTi(ALUDSTRegA), .A(ALUARegA), .B(ALUBRegA), .C(ALUCRegA), .D(ALUDRegA),
				.OpCODE(ALUOpCODERegA), .SA(ALUSARegA), .SB(ALUSBRegA), .SC(ALUSCRegA), .SD(ALUSDRegA), .R(ALURA), .COUT(ALUCOUTA), 
				.DSTo(ALUDSTA), .SR(ALUSRA), .RDY(ALURDYA), .OVR(ALUOVRA), .Zero(ALUZeroA), .Sign(ALUSignA));
ALU64X16 IntALUB (.CLK(CLK), .ACT(ALUACTRegB), .CIN(1'b0), .DSTi(ALUDSTRegB), .A(ALUARegB), .B(ALUBRegB), .C(ALUCRegB), .D(ALUDRegB),
				.OpCODE(ALUOpCODERegB), .SA(ALUSARegB), .SB(ALUSBRegB), .SC(ALUSCRegB), .SD(ALUSDRegB), .R(ALURB), .COUT(ALUCOUTB),
				.DSTo(ALUDSTB), .SR(ALUSRB), .RDY(ALURDYB), .OVR(ALUOVRB), .Zero(ALUZeroB), .Sign(ALUSignB));

// shifter
Shifter64X16 Sht (.CLK(CLK), .ACT(ShiftACTReg), .CIN(0), .A(ShiftAReg), .B(ShiftBReg), .DSTi(ShiftDSTReg),
				.SA(ShiftSAReg), .OPR(ShiftOPRReg), .R(ShiftR), .DSTo(ShiftDST), .RDY(ShiftRDY), .OVR(ShiftOVR),
				.ZERO(ShiftZERO), .SIGN(ShiftSign), .COUT(ShiftCOUT), .SR(ShiftSR));

// misc unit
Misc64X16 Misc (.CLK(CLK), .ACT(MiscACTReg), .OpCODE(MiscOPRReg), .SA(MiscSAReg), .SD(MiscSDReg), .DSTi(MiscDSTReg),
				.CIN(MiscCINReg), .A(MiscAReg), .RDY(MiscRDY), .ZERO(MiscZero), .NaN(MiscNaN), .SIGN(MiscSign),
				.OVR(MiscOVR), .COUT(MiscCOUT), .SR(MiscSR), .DSTo(MiscDST), .R(MiscR));

/*
===========================================================================================================
				Assignments part
===========================================================================================================
*/
assign RIP={PrefRealIP, 1'b0};

// error reporting
assign ESTB=(((DLMachine==ZSS) | (DLMachine==INVSS) | (DLMachine==AERSS)) & ~CheckTag[6] & ~CheckTag[5]) | CodeError | (DLMachine==INVOBS);
assign ECD[23:0]=CodeError ? ADR[13][23:0] : ((DLMachine==INVOBS) ? InvalidSelector : CheckSelector[23:0]);
assign ECD[24]=CodeError | LoadLowerDSC | LoadUpperDSC;
assign ECD[25]=CodeError | (DLMachine==AERSS);
assign ECD[26]=InvalidCPL & ~CodeError;
assign ECD[27]=InvalidTaskID & ~CodeError;
assign ECD[28]=InvalidType & ~CodeError;

assign CSEL=ADR[13][23:0];

/*
===========================================================================================================
				Asynchronous part
===========================================================================================================
*/
always @*
	begin
	
	// LOOP instruction flag
	LoopInstFlag=MiscInstReg[3] & MiscInstReg[2] & MiscInstReg[1] & MiscInstReg[0];

	// Next node on the check access stage
	CheckNext=(~ACT | NEXT) & (~StreamACT | StreamNEXT) & (~NetACT | NetNEXT);
	
	// next node on the memory forming stage
	MemNext=~CheckACT | (CheckNext & ((CheckAR[3] & (CheckOffset[36:5]>=CheckLL) & (CheckOffset[36:5]<CheckUL) & (CheckCMD | CheckAR[1]) & 
													(~CheckCMD | CheckAR[0])) | (CheckAR[3] & CheckAR[2]) | CheckNetwork)) |
						((DLMachine==STS) & (~CheckTag[6] | ~CheckTag[5] | CheckTag[4] | CheckTag[3] | CheckNext));
	
	// forming condition code for prefetcher
	case (PrefInstReg[11:9])
		3'd0:	PrefCC=PrefInstReg[12] ^ ((AFR[PrefInstReg[8:5]][16] & ~(|PrefCCBypassReg)) | (FADDZeroA & PrefCCBypassReg[0]) | (FMULZeroA[0] & PrefCCBypassReg[1]) |
										(FMULZeroA[1] & PrefCCBypassReg[2]) | (ALUZeroA & PrefCCBypassReg[3]) | (ShiftZERO & PrefCCBypassReg[4]) | (MiscZero & PrefCCBypassReg[5]) |
										(FADDZeroB & PrefCCBypassReg[6]) | (FMULZeroB[0] & PrefCCBypassReg[7]) | (FMULZeroB[1] & PrefCCBypassReg[8]) |
										(ALUZeroB & PrefCCBypassReg[9]));
		3'd1:	PrefCC=PrefInstReg[12] ^ ((AFR[PrefInstReg[8:5]][15] & ~PrefCCBypassReg[3] & ~PrefCCBypassReg[5] & ~PrefCCBypassReg[9]) |
										(ALUCOUTA[15] & PrefCCBypassReg[3]) | (MiscCOUT & PrefCCBypassReg[5]) | (ALUCOUTB[15] & PrefCCBypassReg[9]));
		3'd2:	PrefCC=PrefInstReg[12] ^ ((AFR[PrefInstReg[8:5]][17] & ~(|PrefCCBypassReg)) | (FADDSignA & PrefCCBypassReg[0]) | (FMULSignA[0] & PrefCCBypassReg[1]) |
										(FMULSignA[1] & PrefCCBypassReg[2]) | (ALUSignA & PrefCCBypassReg[3]) | (ShiftSign & PrefCCBypassReg[4]) | (MiscSign & PrefCCBypassReg[5]) |
										(FADDSignB & PrefCCBypassReg[6]) | (FMULSignB[0] & PrefCCBypassReg[7]) | (FMULSignB[1] & PrefCCBypassReg[8]) | (ALUSignB & PrefCCBypassReg[9]));
		3'd3:	PrefCC=PrefInstReg[12] ^ ((AFR[PrefInstReg[8:5]][18] & ~PrefCCBypassReg[3] & ~PrefCCBypassReg[4] & ~PrefCCBypassReg[9]) |
										(ALUOVRA & PrefCCBypassReg[3]) | (ShiftOVR & PrefCCBypassReg[4]) | (ALUOVRB & PrefCCBypassReg[9]));
		3'd4:	PrefCC=PrefInstReg[12] ^ ((AFR[PrefInstReg[8:5]][19] & ~PrefCCBypassReg[0] & ~PrefCCBypassReg[1] & ~PrefCCBypassReg[2] & ~PrefCCBypassReg[5] &
										~PrefCCBypassReg[6] & ~PrefCCBypassReg[7] & ~PrefCCBypassReg[8]) |
										(FADDInfA & PrefCCBypassReg[0]) | (FMULInfA[0] & PrefCCBypassReg[1]) | (FMULInfA[1] & PrefCCBypassReg[2]) | (MiscOVR & PrefCCBypassReg[5]) |
										(FADDInfB & PrefCCBypassReg[6]) | (FMULInfB[0] & PrefCCBypassReg[7]) | (FMULInfB[1] & PrefCCBypassReg[8]));
		3'd5:	PrefCC=PrefInstReg[12] ^ ((AFR[PrefInstReg[8:5]][20] & ~PrefCCBypassReg[0] & ~PrefCCBypassReg[1] & ~PrefCCBypassReg[2] & ~PrefCCBypassReg[5] &
										~PrefCCBypassReg[6] & ~PrefCCBypassReg[7] & ~PrefCCBypassReg[8]) |
										(FADDNaNA & PrefCCBypassReg[0]) | (FMULNaNA[0] & PrefCCBypassReg[1]) | (FMULNaNA[1] & PrefCCBypassReg[2]) | (MiscNaN & PrefCCBypassReg[5]) |
										(FADDNaNB & PrefCCBypassReg[6]) | (FMULNaNB[0] & PrefCCBypassReg[7]) | (FMULNaNB[1] & PrefCCBypassReg[8]));
		3'd6:	PrefCC=PrefInstReg[12] ^ ((AFR[PrefInstReg[8:5]][21] & ~PrefCCBypassReg[4]) | (ShiftCOUT & PrefCCBypassReg[4]));
		3'd7:	PrefCC=1'b1;
		endcase

	// forming flags for reset LI counters
	for (i=0; i<16; i=i+1)
		LIResetFlag[i]=(FADDInstRegA[0] & ((FADDInstRegA[5:2]==i) | (FADDInstRegA[9:6]==i) | (FADDInstRegA[13:10]==i)))|
						(FADDInstRegB[0] & ((FADDInstRegB[5:2]==i) | (FADDInstRegB[9:6]==i) | (FADDInstRegB[13:10]==i)))|
						(FMULInstRegA[0] & ((FMULInstRegA[4:1]==i) | (FMULInstRegA[8:5]==i) | (FMULInstRegA[12:9]==i)))|
						(FMULInstRegB[0] & ((FMULInstRegB[4:1]==i) | (FMULInstRegB[8:5]==i) | (FMULInstRegB[12:9]==i)))|
						(FMULACCReg[0] & ((FMULACCReg[7:4]==i) | (FMULACCReg[11:8]==i) | (FMULACCReg[15:12]==i)))|
						(FDIVInstReg[0] & (((FDIVInstReg[4:1]==i) & ~FDIVInstReg[13]) | (FDIVInstReg[8:5]==i) | (FDIVInstReg[12:9]==i)))|
						(ALUInstRegA[0] & (((ALUInstRegA[6:3]==i) & ~ALUInstRegA[15]) | ((ALUInstRegA[10:7]==i) & ~ALUInstRegA[15]) | 
											((ALUInstRegA[14:11]==i) & ~ALUInstRegA[24]) | ((ALUInstRegA[23:20]==i) & ALUInstRegA[24]) |
											((ALUInstRegA[19:16]==i) & ALUInstRegA[24])))|
						(ALUInstRegB[0] & (((ALUInstRegB[6:3]==i) & ~ALUInstRegB[15]) | ((ALUInstRegB[10:7]==i) & ~ALUInstRegB[15]) | 
											((ALUInstRegB[14:11]==i) & ~ALUInstRegB[24]) | ((ALUInstRegB[23:20]==i) & ALUInstRegB[24]) |
											((ALUInstRegB[19:16]==i) & ALUInstRegB[24])))|
						(ShiftInstReg[0] & ((ShiftInstReg[12:9]==i) | (ShiftInstReg[4] & (ShiftInstReg[8:5]==i))))|
						(MiscInstReg[0] & ((MiscInstReg[11:8]==i) | (MiscInstReg[3] & ~(MiscInstReg[2] & MiscInstReg[1]) & (MiscInstReg[7:4]==i))))|
						(MovInstReg[0] & (((MovInstReg[14:11]==i) & (MovInstReg[2:1]!=2'b11)) | ((MovInstReg[10:7]==i) & (MovInstReg[2:1]==2'b00))))|
						(PrefInstReg[0] & (((PrefInstReg[8:5]==i) & (PrefInstReg[4:1]==4'd2)) | 
											((PrefInstReg[16:13]==i) & (PrefInstReg[8:1]==8'hF0) & 
																	((PrefInstReg[12:10]==3'd3) | (PrefInstReg[12:10]==3'd5) | (PrefInstReg[12:9]==4'hC)))))|
						(MemInstReg[0] & (((MemInstReg[15:12]==i) & (MemInstReg[4:1]!=4'd6) & (~(MemInstReg[11] & (&MemInstReg[3:1])))) | 
											((MemInstReg[11:8]==i) & ((MemInstReg[4:3]==2'b10) | 
																														(MemInstReg[4:1]==4'b1100) |
																														(MemInstReg[4:1]==4'b0000) |
																														(MemInstReg[4:1]==4'b0110)))));

	// Memory operand Size forming
	MemoryOSValue[4]=MemLDST & (MemSize==3'b100);
	MemoryOSValue[3]=MemPUSH | MemPOP | (MemLDST & (MemSize==3'b011));
	MemoryOSValue[2]=MemLDST & (MemSize==3'b010);
	MemoryOSValue[1]=MemLDST & (MemSize==3'b001);
	MemoryOSValue[0]=MemLDST & (MemSize==3'b000);

	// interface to the descriptor reloading system
	// Load New sel flag
	LoadNewDSC=CheckACT & ~CheckAR[3] & ~CheckNetwork;
	// load lower segment
	LoadLowerDSC=CheckACT & CheckAR[3] & ~CheckAR[2] & (CheckOffset[36:5]<CheckLL) & ~CheckNetwork;
	// load upper segment
	LoadUpperDSC=CheckACT & CheckAR[3] & ~CheckAR[2] & (CheckOffset[36:5]>=CheckUL) & ~CheckNetwork;
	// access error by type
	AccessError=CheckACT & CheckAR[3] & ~CheckNetwork & ((~CheckCMD & ~CheckAR[1]) | (CheckCMD & ~CheckAR[0])) & ~CheckPref;

	end

/*
===========================================================================================================
				Synchronous part
===========================================================================================================
*/
always @(negedge RESET or posedge CLK)
if (!RESET) begin
				LIFlag<=16'd0;
				GPVFReg<=16'hFFFF;
				AFR[0]<=32'd0;
				AFR[1]<=32'd0;
				AFR[2]<=32'd0;
				AFR[3]<=32'd0;
				AFR[4]<=32'd0;
				AFR[5]<=32'd0;
				AFR[6]<=32'd0;
				AFR[7]<=32'd0;
				AFR[8]<=32'd0;
				AFR[9]<=32'd0;
				AFR[10]<=32'd0;
				AFR[11]<=32'd0;
				AFR[12]<=32'd0;
				AFR[13]<=32'd0;
				AFR[14]<=32'd0;
				AFR[15]<=32'd0;
				ADR[0]<=0;
				ADR[1]<=0;
				ADR[2]<=0;
				ADR[3]<=0;
				ADR[4]<=0;
				ADR[5]<=0;
				ADR[6]<=0;
				ADR[7]<=0;
				ADR[8]<=0;
				ADR[9]<=0;
				ADR[10]<=0;
				ADR[11]<=0;
				ADR[12]<=0;
				ADR[13]<=0;
				ADR[14]<=0;
				ADR[15]<=0;
				GPR[0]<=0;
				GPR[1]<=0;
				GPR[2]<=0;
				GPR[3]<=0;
				GPR[4]<=0;
				GPR[5]<=0;
				GPR[6]<=0;
				GPR[7]<=0;
				GPR[8]<=0;
				GPR[9]<=0;
				GPR[10]<=0;
				GPR[11]<=0;
				GPR[12]<=0;
				GPR[13]<=0;
				GPR[14]<=0;
				GPR[15]<=0;
				FMULACCReg[0]<=1'b0;
				FADDInstRegA[0]<=1'b0;
				FADDInstRegB[0]<=1'b0;
				FMULInstRegA[0]<=1'b0;
				FMULInstRegB[0]<=1'b0;
				FDIVInstReg[0]<=1'b0;
				FDIVACTReg<=1'b0;
				ALUInstRegA[0]<=1'b0;
				ALUInstRegB[0]<=1'b0;
				ShiftInstReg[0]<=1'b0;
				MiscInstReg[0]<=1'b0;
				LoopInstReg[0]<=1'b0;
				PrefInstReg[0]<=1'b0;
				MovInstReg[0]<=1'b0;
				MemInstReg[0]<=1'b0;
				MemBusy<=1'b0;
				MemCNT<=2'b00;
				CheckACT<=1'b0;
				ACT<=1'b0;
				StreamACT<=1'b0;
				NetACT<=1'b0;
				DLMachine<=WS;
				DescriptorLoadState<=1'b0;
				DTR[0]<=156'hB000000000000FFFFFFFF000000000000000000;
				DTR[1]<=156'hB000000000000FFFFFFFF000000000000000000;
				DTR[2]<=156'hB000000000000FFFFFFFF000000000000000000;
				DTR[3]<=156'hB000000000000FFFFFFFF000000000000000000;
				DTR[4]<=156'hB000000000000FFFFFFFF000000000000000000;
				DTR[5]<=156'hB000000000000FFFFFFFF00000000FFFFFFFFFC;
				DTR[6]<=156'hB000000000000FFFFFFFF000000000000000000;
				DTR[7]<=156'hB000000000000FFFFFFFF000000000000000000;
				PrefCallReg<=1'b0;
				PrefRetReg<=1'b0;
				MemReadAR<=0;
				MemLoadOffset<=0;
				MemLoadSel<=0;
				MemReq<=0;
				MemPUSH<=0;
				MemPOP<=0;
				MemADRPushPop<=0;
				MemLDO<=0;
				FMULACCACTReg<=0;
				FMULACCDRDYFlag<=0;
				FFT32NEXTReg<=0;
				IV<=0;
				MemFifoFullFlag<=0;
				end
else begin
	
	// Fifo full flag
	MemFifoFullFlag<=(MemFifoUsedW>6'd59);
	
	// Instructions transfered to the sequencer
	IV<=IVF & {4{IFetch & InsRDY}};

	// EU empty flag
	EMPTY<=PrefEMPTY & SeqEMPTY & (&GPVFReg);
	
	// output data for context store operations
	case (RA[5:4])
		2'd0: CDATA<=GPR[RA[3:0]][63:0];
		2'd1: CDATA<=GPR[RA[3:0]][127:64];
		2'd2: CDATA<={32'd0, AFR[RA[3:0]]};
		2'd3: CDATA<={27'd0, ADR[RA[3:0]]};
		endcase
	
	// Storing TAGi
	TAGiReg<=TAGi;

	// LI flags
	for (i=0; i<16; i=i+1)
		LIFlag[i]<=(&MovInstReg[2:0]) & (MovInstReg[14:11]==i);
	
	// processign GPR valid flags
	for (i=0; i<16; i=i+1)
			GPVFReg[i]<=(GPVFReg[i] & GPVFINVD[i])|
						((FADDDSTA==i) & FADDRDYA)|
						((FADDDSTB==i) & FADDRDYB)|
						((FMULDSTA[0]==i) & FMULRDYA[0])|
						((FMULDSTA[1]==i) & FMULRDYA[1])|
						((FMULDSTB[0]==i) & FMULRDYB[0])|
						((FMULDSTB[1]==i) & FMULRDYB[1])|
						FMULACCSelNode[i]|
						((FMULACCDSTReg==i) & FMULACCACTReg & FMULACCCMDReg)|
						((FDIVDST==i) & FDIVRDY)|
						((ALUDSTA==i) & ALURDYA)|
						((ALUDSTB==i) & ALURDYB)|
						((ShiftDST==i) & ShiftRDY)|
						((MiscDST==i) & MiscRDY)|
						((MovInstReg[14:11]==i) & MovInstReg[0])|
						(MemReadAR & (MemDST==i))|
						(DRDY & (TAGi[3:0]==i) & ~TAGi[6] & ~TAGi[5] & (~TAGi[7] | TAGi[4])) |
						(SkipDataRead & (STAGReg==i));
	// result strobe nodes
	for (i=0; i<16; i=i+1)
		begin
		FlagWrite[i]<=(FADDRDYRA & (FADDDSTRA==i))|
						(FADDRDYRB & (FADDDSTRB==i))|
						(FMULRDYRA[0] & (FMULDSTRA[0]==i))|
						(FMULRDYRA[1] & (FMULDSTRA[1]==i))|
						(FMULRDYRB[0] & (FMULDSTRB[0]==i))|
						(FMULRDYRB[1] & (FMULDSTRB[1]==i))|
						(FMULACCRDY & (FMULACCDST==i))|
						(FMULACCACTReg & FMULACCCMDReg & (FMULACCDSTReg==i))|
						(FDIVRDY & (FDIVDST==i))|
						(ALURDYRA & (ALUDSTRA==i))|
						(ALURDYRB & (ALUDSTRB==i))|
						(ShiftRDYR & (ShiftDSTR==i))|
						(MiscRDYR & (MiscDSTR==i))|
						(DRDY & (TAGi[3:0]==i) & ~TAGi[6] & ((TAGi[5] & ~TAGi[4]) | (~TAGi[5] & (~TAGi[7] | TAGi[4]))));

		GPRByteNode[i]<=(FADDRDYRA & (FADDDSTRA==i))|
						(FADDRDYRB & (FADDDSTRB==i))|
						(FMULRDYRA[0] & (FMULDSTRA[0]==i))|
						(FMULRDYRA[1] & (FMULDSTRA[1]==i))|
						(FMULRDYRB[0] & (FMULDSTRB[0]==i))|
						(FMULRDYRB[1] & (FMULDSTRB[1]==i))|
						(FMULACCRDY & (FMULACCDST==i))|
						(FDIVRDY & (FDIVDST==i))|
						(ALURDYRA & (ALUDSTRA==i))|
						(ALURDYRB & (ALUDSTRB==i))|
						(ShiftRDYR & (ShiftDSTR==i))|
						(MiscRDYR & (MiscDSTR==i))|
						(MovInstReg[0] & (MovInstReg[14:11]==i) & (MovInstReg[2:1]!=2'b01))|
						(MemReadAR & (MemDST==i))|
						(DRDY & (TAGi[3:0]==i) & ~TAGi[6] & ~TAGi[5] & ~TAGi[4]);

		GPRWordNode[i]<=(FADDRDYRA & (FADDDSTRA==i))|
						(FADDRDYRB & (FADDDSTRB==i))|
						(FMULRDYRA[0] & (FMULDSTRA[0]==i))|
						(FMULRDYRA[1] & (FMULDSTRA[1]==i))|
						(FMULRDYRB[0] & (FMULDSTRB[0]==i))|
						(FMULRDYRB[1] & (FMULDSTRB[1]==i))|
						(FMULACCRDY & (FMULACCDST==i))|
						(FDIVRDY & (FDIVDST==i))|
						(ALURDYRA & (ALUDSTRA==i) & (|ALUSRA))|
						(ALURDYRB & (ALUDSTRB==i) & (|ALUSRB))|
						(ShiftRDYR & (ShiftDSTR==i) & (|ShiftSR))|
						(MiscRDYR & (MiscDSTR==i) & (|MiscSR))|
						(MovInstReg[0] & (MovInstReg[14:11]==i) & (MovInstReg[2:1]!=2'b01))|
						(MemReadAR & (MemDST==i))|
						(DRDY & (TAGi[3:0]==i) & (|SZi[1:0]) & ~TAGi[6] & ~TAGi[5] & ~TAGi[4]);

		GPRDwordNode[i]<=(FADDRDYRA & (FADDDSTRA==i))|
						(FADDRDYRB & (FADDDSTRB==i))|
						(FMULRDYRA[0] & (FMULDSTRA[0]==i))|
						(FMULRDYRA[1] & (FMULDSTRA[1]==i))|
						(FMULRDYRB[0] & (FMULDSTRB[0]==i))|
						(FMULRDYRB[1] & (FMULDSTRB[1]==i))|
						(FMULACCRDY & (FMULACCDST==i))|
						(FDIVRDY & (FDIVDST==i))|
						(ALURDYRA & (ALUDSTRA==i) & ALUSRA[1])|
						(ALURDYRB & (ALUDSTRB==i) & ALUSRB[1])|
						(ShiftRDYR & (ShiftDSTR==i) & ShiftSR[1])|
						(MiscRDYR & (MiscDSTR==i) & (MiscSR[2] | MiscSR[1]))|
						(MovInstReg[0] & (MovInstReg[14:11]==i) & (MovInstReg[2:1]!=2'b01))|
						(MemReadAR & (MemDST==i))|
						(DRDY & (TAGi[3:0]==i)& SZi[1] & ~TAGi[6] & ~TAGi[5] & ~TAGi[4]);

		GPRQwordNode[i]<=(FADDRDYRA & (FADDDSTRA==i))|
						(FADDRDYRB & (FADDDSTRB==i))|
						(FMULRDYRA[0] & (FMULDSTRA[0]==i))|
						(FMULRDYRA[1] & (FMULDSTRA[1]==i))|
						(FMULRDYRB[0] & (FMULDSTRB[0]==i))|
						(FMULRDYRB[1] & (FMULDSTRB[1]==i))|
						(FDIVRDY & (FDIVDST==i) & (FDIVSR[2] | FDIVSR[0]))|
						(ALURDYRA & (ALUDSTRA==i) & (&ALUSRA))|
						(ALURDYRB & (ALUDSTRB==i) & (&ALUSRB))|
						(ShiftRDYR & (ShiftDSTR==i) & ShiftSR[1] & ShiftSR[0])|
						(MiscRDYR & (MiscDSTR==i) & ((MiscSR[1] & MiscSR[0]) | MiscSR[2]))|
						(MovInstReg[0] & (MovInstReg[14:11]==i) & (MovInstReg[2:1]!=2'b01))|
						(MemReadAR & (MemDST==i))|
						(DRDY & (TAGi[3:0]==i) & (&SZi[1:0]) & ~TAGi[6] & ~TAGi[5] & ~TAGi[4]);
		
		GPROwordNode[i]<=(MovInstReg[0] & (MovInstReg[14:11]==i) & (MovInstReg[2:1]!=2'b01))|
						(FMULRDYRA[1] & (FMULDSTRA[1]==i))|
						(FMULRDYRB[1] & (FMULDSTRB[1]==i))|
						(FDIVRDY & (FDIVDST==i) & FDIVSR[2])|
						(FADDRDYRA & (FADDDSTRA==i))|
						(FADDRDYRB & (FADDDSTRB==i))|
						(MiscRDYR & (MiscDSTR==i) & MiscSR[2])|
						(DRDY & (TAGi[3:0]==i) & ~TAGi[6] & ~TAGi[5] & TAGi[4]);
		end
	// data selection nodes
	for (i=0; i<16; i=i+1)
		begin
		FADDSelNodeA[i]<=FADDRDYRA & (FADDDSTRA==i);
		FADDSelNodeB[i]<=FADDRDYRB & (FADDDSTRB==i);
		FMULSelNodeA[i]<=FMULRDYRA[0] & (FMULDSTRA[0]==i);
		FMULQSelNodeA[i]<=FMULRDYRA[1] & (FMULDSTRA[1]==i);
		FMULSelNodeB[i]<=FMULRDYRB[0] & (FMULDSTRB[0]==i);
		FMULQSelNodeB[i]<=FMULRDYRB[1] & (FMULDSTRB[1]==i);
		FMULACCSelNode[i]<=FMULACCRDY & (FMULACCDST==i);
		FFTSelNode[i]<=FMULACCACTReg & FMULACCCMDReg & (FMULACCDSTReg==i);
		FDIVSelNode[i]<=FDIVRDY & (FDIVDST==i);
		ALUSelNodeA[i]<=ALURDYRA & (ALUDSTRA==i);
		ALUSelNodeB[i]<=ALURDYRB & (ALUDSTRB==i);
		ShiftSelNode[i]<=ShiftRDYR & (ShiftDSTR==i);
		MiscSelNode[i]<=MiscRDYR & (MiscDSTR==i);
		MovSelNode[i]<=(MovInstReg[0] & (MovInstReg[14:11]==i) & (MovInstReg[2:1]!=2'b01));
		MemSelNode[i]<=DRDY & (TAGi[3:0]==i) & ~TAGi[6] & ~TAGi[5];
		MemFSelNode[i]<=DRDY & (TAGi[3:0]==i) & ~TAGi[6] & TAGi[5] & ~TAGi[4];
		MemASelNode[i]<=DRDY & (TAGi[3:0]==i) & ~TAGi[6] & TAGi[5] & TAGi[4];
		MemARSelNode[i]<=MemReadAR & (MemDST==i);
		end
	// load selector from memory node
	MemLSelNode<=DRDY & ~TAGi[6] & TAGi[0] & TAGi[5] & TAGi[4];

	// DTR selection nodes
	for (i=0; i<8; i=i+1) DTRWriteFlag[i]<=DRDY & ~TAGi[7] & TAGi[6] & ~TAGi[5] &(TAGi[4:2]==i);
	DTRWriteFlag[8]<=DRDY & ~TAGi[7] & TAGi[6] & ~TAGi[5];
	
	// Context loading Flag
	ContextLoadFlag<=CLOAD;	

	// delayed ready registers
	FADDRDYRA<=FADDRDYA;
	FADDRDYRB<=FADDRDYB;
	FMULRDYRA[0]<=FMULRDYA[0];
	FMULRDYRB[0]<=FMULRDYB[0];
	FMULRDYRA[1]<=FMULRDYA[1];
	FMULRDYRB[1]<=FMULRDYB[1];
	ALURDYRA<=ALURDYA;
	ALURDYRB<=ALURDYB;
	ShiftRDYR<=ShiftRDY;
	MiscRDYR<=MiscRDY;
	// delayed destination registers
	FADDDSTRA<=FADDDSTA;
	FADDDSTRB<=FADDDSTB;
	FMULDSTRA[0]<=FMULDSTA[0];
	FMULDSTRB[0]<=FMULDSTB[0];
	FMULDSTRA[1]<=FMULDSTA[1];
	FMULDSTRB[1]<=FMULDSTB[1];
	ALUDSTRA<=ALUDSTA;
	ALUDSTRB<=ALUDSTB;
	ShiftDSTR<=ShiftDST;
	MiscDSTR<=MiscDST;
	// delayed size registers
	FDIVSRReg<=FDIVSR;
	ALUSRRegA<=ALUSRA;
	ALUSRRegB<=ALUSRB;
	ShiftSRReg<=ShiftSR;
	MiscSRReg<=MiscSR;
	SZiReg<=SZi;

	// storing results into registers
	for (i=0; i<16; i=i+1)
		begin
		// storing arithmetic flags
		if (FlagWrite[i])
			begin
			// CF[15:0]
			AFR[i][14:0]<=(ALUCOUTA[14:0] & {15{ALUSelNodeA[i]}}) | (ALUCOUTB[14:0] & {15{ALUSelNodeB[i]}}) | (DTi[14:0] & {15{MemFSelNode[i]}});
			AFR[i][15]<=(ALUCOUTA[15] & ALUSelNodeA[i])|(ALUCOUTB[15] & ALUSelNodeB[i])|(MiscCOUT & MiscSelNode[i])|(DTi[15] & MemFSelNode[i]);
			// ZF
			AFR[i][16]<=(FADDZeroA & FADDSelNodeA[i])|(FADDZeroB & FADDSelNodeB[i])|
						(FMULZeroA[0] & FMULSelNodeA[i])|(FMULZeroA[1] & FMULQSelNodeA[i])|
						(FMULZeroB[0] & FMULSelNodeB[i])|(FMULZeroB[1] & FMULQSelNodeB[i])|
						(FMULACCZERO & FMULACCSelNode[i])|
						(FDIVZero & FDIVSelNode[i])|
						(ALUZeroA & ALUSelNodeA[i])|(ALUZeroB & ALUSelNodeB[i])|
						(ShiftZERO & ShiftSelNode[i])|(MiscZero & MiscSelNode[i])|(DTi[16] & MemFSelNode[i])|
						(FFT32NEXTReg & FFTSelNode[i]);
			// SF
			AFR[i][17]<=(FADDSignA & FADDSelNodeA[i])|(FADDSignB & FADDSelNodeB[i])|
						(FMULSignA[0] & FMULSelNodeA[i])|(FMULSignA[1] & FMULQSelNodeA[i])|
						(FMULSignB[0] & FMULSelNodeB[i])|(FMULSignB[1] & FMULQSelNodeB[i])|
						(FMULACCSIGN & FMULACCSelNode[i])|
						(FDIVSign & FDIVSelNode[i])|
						(ALUSignA & ALUSelNodeA[i])|(ALUSignB & ALUSelNodeB[i])|
						(ShiftSign & ShiftSelNode[i])|(MiscSign & MiscSelNode[i])|(DTi[17] & MemFSelNode[i]);
			// OF
			AFR[i][18]<=(ALUOVRA & ALUSelNodeA[i])|(ALUOVRB & ALUSelNodeB[i])|(ShiftOVR & ShiftSelNode[i])|(DTi[18] & MemFSelNode[i]);
			// IF
			AFR[i][19]<=(FADDInfA & FADDSelNodeA[i])|(FADDInfB & FADDSelNodeB[i])|
						(FMULInfA[0] & FMULSelNodeA[i])|(FMULInfA[1] & FMULQSelNodeA[i])|
						(FMULInfB[0] & FMULSelNodeB[i])|(FMULInfB[1] & FMULQSelNodeB[i])|
						(FMULACCINF & FMULACCSelNode[i])|(FDIVInf & FDIVSelNode[i])|
						(MiscOVR & MiscSelNode[i])|(DTi[19] & MemFSelNode[i]);
			// NF
			AFR[i][20]<=(FADDNaNA & FADDSelNodeA[i])|(FADDNaNB & FADDSelNodeB[i])|
						(FMULNaNA[0] & FMULSelNodeA[i])|(FMULNaNA[1] & FMULQSelNodeA[i])|
						(FMULNaNB[0] & FMULSelNodeB[i])|(FMULNaNB[1] & FMULQSelNodeB[i])|
						(FDIVNaN & FDIVSelNode[i])|(MiscNaN & MiscSelNode[i])|
						(DTi[20] & MemFSelNode[i])|(MemSelNode[i] & (&SZiReg))|
						(FMULACCNAN & FMULACCSelNode[i]);
			// DBF
			AFR[i][21]<=(ShiftCOUT & ShiftSelNode[i])|(DTi[21] & MemFSelNode[i]);
			end
		// Size of operand and address mode
		if (MemFSelNode[i]) AFR[i][27:22]<=DTi[27:22];
			else if (MemSelNode[i]) AFR[i][24:22]<=TAGiReg[7] ? 3'd4 : {SZiReg};
				else if (MovSelNode[i]) AFR[i][24:22]<=MovSR;
					else if (MemARSelNode[i]) AFR[i][24:22]<=3'b011;
						else if (FADDSelNodeA[i] | FADDSelNodeB[i] | FMULSelNodeA[i] | FMULQSelNodeA[i] | FMULSelNodeB[i] | FMULQSelNodeB[i] | FDIVSelNode[i] | ALUSelNodeA[i] | ALUSelNodeB[i] | ShiftSelNode[i] | MiscSelNode[i] | FMULACCSelNode[i])
							begin
							AFR[i][24]<=FMULQSelNodeA[i] | FMULQSelNodeB[i] | (FADDSRA[2] & FADDSelNodeA[i]) | (FADDSRB[2] & FADDSelNodeB[i]) | (MiscSRReg[2] & MiscSelNode[i]) | (FDIVSRReg[2] & FDIVSelNode[i]);
							AFR[i][23:22]<=(FADDSRA[1:0] & {2{FADDSelNodeA[i]}})|
										(FADDSRB[1:0] & {2{FADDSelNodeB[i]}})|
										({1'b1, FMULSRA} & {2{FMULSelNodeA[i]}})|
										({1'b1, FMULSRB} & {2{FMULSelNodeB[i]}})|
										(FDIVSRReg[1:0] & {2{FDIVSelNode[i]}})|
										(ALUSRRegA & {2{ALUSelNodeA[i]}})|
										(ALUSRRegB & {2{ALUSelNodeB[i]}})|
										(ShiftSRReg & {2{ShiftSelNode[i]}})|
										(MiscSRReg[1:0] & {2{MiscSelNode[i]}})| {FMULACCSelNode[i], 1'b0};
							end
		//LI byte counter
		if (LIResetFlag[i] | LIRESET) AFR[i][31:28]<=4'b0000;
			else if (MemFSelNode[i]) AFR[i][31:28]<=DTi[31:28] & {4{ContextLoadFlag}};
				else if (LIFlag[i]) AFR[i][31:28]<=AFR[i][31:28]+4'd1;

		// GPR Bits 7:0
		if (GPRByteNode[i]) GPR[i][7:0]<=(FADDRA[7:0] & {8{FADDSelNodeA[i]}})|
											(FADDRB[7:0] & {8{FADDSelNodeB[i]}})|
											(FMULRA[7:0] & {8{FMULSelNodeA[i]}})|
											(FMULRQA[7:0] & {8{FMULQSelNodeA[i]}})|
											(FMULRB[7:0] & {8{FMULSelNodeB[i]}})|
											(FMULRQB[7:0] & {8{FMULQSelNodeB[i]}})|
											(FMULACCR[7:0] & {8{FMULACCSelNode[i]}})|
											(FDIVR[7:0] & {8{FDIVSelNode[i]}})|
											(ALURA[7:0] & {8{ALUSelNodeA[i]}})|
											(ALURB[7:0] & {8{ALUSelNodeB[i]}})|
											(ShiftR[7:0] & {8{ShiftSelNode[i]}})|
											(MiscR[7:0] & {8{MiscSelNode[i]}})|
											(MovReg[7:0] & {8{MovSelNode[i]}})|
											(DTi[7:0] & {8{MemSelNode[i]}})|
											(ARData[7:0] & {8{MemARSelNode[i]}});
		// GPR Bits 15:8
		if (GPRWordNode[i]) GPR[i][15:8]<=(FADDRA[15:8] & {8{FADDSelNodeA[i]}})|
											(FADDRB[15:8] & {8{FADDSelNodeB[i]}})|
											(FMULRA[15:8] & {8{FMULSelNodeA[i]}})|
											(FMULRQA[15:8] & {8{FMULQSelNodeA[i]}})|
											(FMULRB[15:8] & {8{FMULSelNodeB[i]}})|
											(FMULRQB[15:8] & {8{FMULQSelNodeB[i]}})|
											(FMULACCR[15:8] & {8{FMULACCSelNode[i]}})|
											(FDIVR[15:8] & {8{FDIVSelNode[i]}})|
											(ALURA[15:8] & {8{ALUSelNodeA[i]}})|
											(ALURB[15:8] & {8{ALUSelNodeB[i]}})|
											(ShiftR[15:8] & {8{ShiftSelNode[i]}})|
											(MiscR[15:8] & {8{MiscSelNode[i]}})|
											(MovReg[15:8] & {8{MovSelNode[i]}})|
											(DTi[15:8] & {8{MemSelNode[i]}})|
											(ARData[15:8] & {8{MemARSelNode[i]}});

		if (GPRDwordNode[i]) GPR[i][31:16]<=(FADDRA[31:16] & {16{FADDSelNodeA[i]}})|
											(FADDRB[31:16] & {16{FADDSelNodeB[i]}})|
											(FMULRA[31:16] & {16{FMULSelNodeA[i]}})|
											(FMULRQA[31:16] & {16{FMULQSelNodeA[i]}})|
											(FMULRB[31:16] & {16{FMULSelNodeB[i]}})|
											(FMULRQB[31:16] & {16{FMULQSelNodeB[i]}})|
											(FMULACCR[31:16] & {16{FMULACCSelNode[i]}})|
											(FDIVR[31:16] & {16{FDIVSelNode[i]}})|
											(ALURA[31:16] & {16{ALUSelNodeA[i]}})|
											(ALURB[31:16] & {16{ALUSelNodeB[i]}})|
											(ShiftR[31:16] & {16{ShiftSelNode[i]}})|
											(MiscR[31:16] & {16{MiscSelNode[i]}})|
											(MovReg[31:16] & {16{MovSelNode[i]}})|
											(DTi[31:16] & {16{MemSelNode[i]}})|
											(ARData[31:16] & {16{MemARSelNode[i]}});

		if (GPRQwordNode[i]) GPR[i][63:32]<=(FADDRA[63:32] & {32{FADDSelNodeA[i]}})|
											(FADDRB[63:32] & {32{FADDSelNodeB[i]}})|
											(FMULRA[63:32] & {32{FMULSelNodeA[i]}})|
											(FMULRQA[63:32] & {32{FMULQSelNodeA[i]}})|
											(FMULRB[63:32] & {32{FMULSelNodeB[i]}})|
											(FMULRQB[63:32] & {32{FMULQSelNodeB[i]}})|
											(FDIVR[63:32] & {32{FDIVSelNode[i]}})|
											(ALURA[63:32] & {32{ALUSelNodeA[i]}})|
											(ALURB[63:32] & {32{ALUSelNodeB[i]}})|
											(ShiftR[63:32] & {32{ShiftSelNode[i]}})|
											(MiscR[63:32] & {32{MiscSelNode[i]}})|
											(MovReg[63:32] & {32{MovSelNode[i]}})|
											(DTi[63:32] & {32{MemSelNode[i]}})|
											(ARData[36:32] & {32{MemARSelNode[i]}});
		
		if (GPROwordNode[i]) GPR[i][127:64]<=(MovReg[127:64] & {64{MovSelNode[i]}})|
											(DTi & {64{MemSelNode[i]}})|
											(FMULRQA[127:64] & {64{FMULQSelNodeA[i]}})|
											(FMULRQB[127:64] & {64{FMULQSelNodeB[i]}})|
											(FDIVR[127:64] & {64{FDIVSelNode[i]}})|
											(FADDRA[127:64] & {64{FADDSelNodeA[i]}}) |
											(FADDRB[127:64] & {64{FADDSelNodeB[i]}}) |
											(MiscR[127:64] & {64{MiscSelNode[i]}});
		end

	// processing source operands
	// FADD Channel
	FADDInstRegA<=FADDInstBusA;
	FADDInstRegB<=FADDInstBusB;
	FADDACTRegA<=FADDInstRegA[0];
	FADDACTRegB<=FADDInstRegB[0];
	FADDCMDRegA<=FADDInstRegA[1];
	FADDCMDRegB<=FADDInstRegB[1];

	FADDBypassARegA[0]<=FADDRDYRA & (FADDDSTRA==FADDInstBusA[5:2]);
	FADDBypassARegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FADDInstBusA[5:2]);
	FADDBypassARegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FADDInstBusA[5:2]);
	FADDBypassARegA[3]<=ALURDYRA & (ALUDSTRA==FADDInstBusA[5:2]);
	FADDBypassARegA[4]<=ShiftRDYR & (ShiftDSTR==FADDInstBusA[5:2]);
	FADDBypassARegA[5]<=MiscRDYR & (MiscDSTR==FADDInstBusA[5:2]);
	FADDBypassARegA[6]<=FADDRDYRB & (FADDDSTRB==FADDInstBusA[5:2]);
	FADDBypassARegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FADDInstBusA[5:2]);
	FADDBypassARegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FADDInstBusA[5:2]);
	FADDBypassARegA[9]<=ALURDYRB & (ALUDSTRB==FADDInstBusA[5:2]);

	FADDBypassARegB[0]<=FADDRDYRA & (FADDDSTRA==FADDInstBusB[5:2]);
	FADDBypassARegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FADDInstBusB[5:2]);
	FADDBypassARegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FADDInstBusB[5:2]);
	FADDBypassARegB[3]<=ALURDYRA & (ALUDSTRA==FADDInstBusB[5:2]);
	FADDBypassARegB[4]<=ShiftRDYR & (ShiftDSTR==FADDInstBusB[5:2]);
	FADDBypassARegB[5]<=MiscRDYR & (MiscDSTR==FADDInstBusB[5:2]);
	FADDBypassARegB[6]<=FADDRDYRB & (FADDDSTRB==FADDInstBusB[5:2]);
	FADDBypassARegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FADDInstBusB[5:2]);
	FADDBypassARegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FADDInstBusB[5:2]);
	FADDBypassARegB[9]<=ALURDYRB & (ALUDSTRB==FADDInstBusB[5:2]);

	FADDARegA<=(GPR[FADDInstRegA[5:2]] & {128{~(|FADDBypassARegA)}}) |
				(FADDRA & {128{FADDBypassARegA[0]}}) |
				({64'd0, FMULRA & {64{FADDBypassARegA[1]}}}) |
				(FMULRQA & {128{FADDBypassARegA[2]}}) |
				({GPR[FADDInstRegA[5:2]][127:64], ALURA} & {128{FADDBypassARegA[3]}}) |
				({GPR[FADDInstRegA[5:2]][127:64], ShiftR} & {128{FADDBypassARegA[4]}}) |
				(MiscR & {128{FADDBypassARegA[5]}}) |
				(FADDRB & {128{FADDBypassARegA[6]}}) |
				({64'd0, FMULRB & {64{FADDBypassARegA[7]}}}) |
				(FMULRQB & {128{FADDBypassARegA[8]}}) |
				({GPR[FADDInstRegA[5:2]][127:64], ALURB} & {128{FADDBypassARegA[9]}});
	
	FADDARegB<=(GPR[FADDInstRegB[5:2]] & {128{~(|FADDBypassARegB)}}) |
				(FADDRA & {128{FADDBypassARegB[0]}}) |
				({64'd0, FMULRA & {64{FADDBypassARegB[1]}}}) |
				(FMULRQA & {128{FADDBypassARegB[2]}}) |
				({GPR[FADDInstRegB[5:2]][127:64], ALURA} & {128{FADDBypassARegB[3]}}) |
				({GPR[FADDInstRegB[5:2]][127:64], ShiftR} & {128{FADDBypassARegB[4]}}) |
				(MiscR & {128{FADDBypassARegB[5]}}) |
				(FADDRB & {128{FADDBypassARegB[6]}}) |
				({64'd0, FMULRB & {64{FADDBypassARegB[7]}}}) |
				(FMULRQB & {128{FADDBypassARegB[8]}}) |
				({GPR[FADDInstRegB[5:2]][127:64], ALURB} & {128{FADDBypassARegB[9]}});
	
	FADDSARegA<=(AFR[FADDInstRegA[5:2]][24:22] & {3{~(|FADDBypassARegA)}}) |
				(FADDSRA & {3{FADDBypassARegA[0]}})|
				({2'd1, FMULSRA} & {3{FADDBypassARegA[1]}})|
				({FADDBypassARegA[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FADDBypassARegA[3]}}})|
				({1'b0, ShiftSRReg & {2{FADDBypassARegA[4]}}})|
				(MiscSRReg & {3{FADDBypassARegA[5]}}) |
				(FADDSRB & {3{FADDBypassARegA[6]}})|
				({2'd1, FMULSRB} & {3{FADDBypassARegA[7]}})|
				({FADDBypassARegA[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FADDBypassARegA[9]}}});

	FADDSARegB<=(AFR[FADDInstRegB[5:2]][24:22] & {3{~(|FADDBypassARegB)}}) |
				(FADDSRA & {3{FADDBypassARegB[0]}})|
				({2'd1, FMULSRA} & {3{FADDBypassARegB[1]}})|
				({FADDBypassARegB[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FADDBypassARegB[3]}}})|
				({1'b0, ShiftSRReg & {2{FADDBypassARegB[4]}}})|
				(MiscSRReg & {3{FADDBypassARegB[5]}}) |
				(FADDSRB & {3{FADDBypassARegB[6]}})|
				({2'd1, FMULSRB} & {3{FADDBypassARegB[7]}})|
				({FADDBypassARegB[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FADDBypassARegB[9]}}});

	FADDBypassBRegA[0]<=FADDRDYRA & (FADDDSTRA==FADDInstBusA[9:6]);
	FADDBypassBRegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FADDInstBusA[9:6]);
	FADDBypassBRegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FADDInstBusA[9:6]);
	FADDBypassBRegA[3]<=ALURDYRA & (ALUDSTRA==FADDInstBusA[9:6]);
	FADDBypassBRegA[4]<=ShiftRDYR & (ShiftDSTR==FADDInstBusA[9:6]);
	FADDBypassBRegA[5]<=MiscRDYR & (MiscDSTR==FADDInstBusA[9:6]);
	FADDBypassBRegA[6]<=FADDRDYRB & (FADDDSTRB==FADDInstBusA[9:6]);
	FADDBypassBRegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FADDInstBusA[9:6]);
	FADDBypassBRegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FADDInstBusA[9:6]);
	FADDBypassBRegA[9]<=ALURDYRB & (ALUDSTRB==FADDInstBusA[9:6]);

	FADDBypassBRegB[0]<=FADDRDYRA & (FADDDSTRA==FADDInstBusB[9:6]);
	FADDBypassBRegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FADDInstBusB[9:6]);
	FADDBypassBRegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FADDInstBusB[9:6]);
	FADDBypassBRegB[3]<=ALURDYRA & (ALUDSTRA==FADDInstBusB[9:6]);
	FADDBypassBRegB[4]<=ShiftRDYR & (ShiftDSTR==FADDInstBusB[9:6]);
	FADDBypassBRegB[5]<=MiscRDYR & (MiscDSTR==FADDInstBusB[9:6]);
	FADDBypassBRegB[6]<=FADDRDYRB & (FADDDSTRB==FADDInstBusB[9:6]);
	FADDBypassBRegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FADDInstBusB[9:6]);
	FADDBypassBRegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FADDInstBusB[9:6]);
	FADDBypassBRegB[9]<=ALURDYRB & (ALUDSTRB==FADDInstBusB[9:6]);

	FADDBRegA<=(GPR[FADDInstRegA[9:6]] & {128{~(|FADDBypassBRegA)}}) |
				(FADDRA & {128{FADDBypassBRegA[0]}}) |
				({64'd0, FMULRA & {64{FADDBypassBRegA[1]}}}) |
				(FMULRQA & {128{FADDBypassBRegA[2]}}) |
				({GPR[FADDInstRegA[9:6]][127:64], ALURA} & {128{FADDBypassBRegA[3]}}) |
				({GPR[FADDInstRegA[9:6]][127:64], ShiftR} & {128{FADDBypassBRegA[4]}}) |
				(MiscR & {128{FADDBypassBRegA[5]}}) |
				(FADDRB & {128{FADDBypassBRegA[6]}}) |
				({64'd0, FMULRB & {64{FADDBypassBRegA[7]}}}) |
				(FMULRQB & {128{FADDBypassBRegA[8]}}) |
				({GPR[FADDInstRegA[9:6]][127:64], ALURB} & {128{FADDBypassBRegA[9]}});	
	
	FADDBRegB<=(GPR[FADDInstRegB[9:6]] & {128{~(|FADDBypassBRegB)}}) |
				(FADDRA & {128{FADDBypassBRegB[0]}}) |
				({64'd0, FMULRA & {64{FADDBypassBRegB[1]}}}) |
				(FMULRQA & {128{FADDBypassBRegB[2]}}) |
				({GPR[FADDInstRegB[9:6]][127:64], ALURA} & {128{FADDBypassBRegB[3]}}) |
				({GPR[FADDInstRegB[9:6]][127:64], ShiftR} & {128{FADDBypassBRegB[4]}}) |
				(MiscR & {128{FADDBypassBRegB[5]}}) |
				(FADDRB & {128{FADDBypassBRegB[6]}}) |
				({64'd0, FMULRB & {64{FADDBypassBRegB[7]}}}) |
				(FMULRQB & {128{FADDBypassBRegB[8]}}) |
				({GPR[FADDInstRegB[9:6]][127:64], ALURB} & {128{FADDBypassBRegB[9]}});

	FADDSBRegA<=(AFR[FADDInstRegA[9:6]][24:22] & {3{~(|FADDBypassBRegA)}})|
				(FADDSRA & {3{FADDBypassBRegA[0]}})|
				({2'd1, FMULSRA} & {3{FADDBypassBRegA[1]}})|
				({FADDBypassBRegA[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FADDBypassBRegA[3]}}})|
				({1'b0, ShiftSRReg & {2{FADDBypassBRegA[4]}}})|
				(MiscSRReg & {3{FADDBypassBRegA[5]}})|
				(FADDSRB & {3{FADDBypassBRegA[6]}})|
				({2'd1, FMULSRB} & {3{FADDBypassBRegA[7]}})|
				({FADDBypassBRegA[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FADDBypassBRegA[9]}}});
	
	FADDSBRegB<=(AFR[FADDInstRegB[9:6]][24:22] & {3{~(|FADDBypassBRegB)}})|
				(FADDSRA & {3{FADDBypassBRegB[0]}})|
				({2'd1, FMULSRA} & {3{FADDBypassBRegB[1]}})|
				({FADDBypassBRegB[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FADDBypassBRegB[3]}}})|
				({1'b0, ShiftSRReg & {2{FADDBypassBRegB[4]}}})|
				(MiscSRReg & {3{FADDBypassBRegB[5]}})|
				(FADDSRB & {3{FADDBypassBRegB[6]}})|
				({2'd1, FMULSRB} & {3{FADDBypassBRegB[7]}})|
				({FADDBypassBRegB[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FADDBypassBRegB[9]}}});
	
	FADDDSTRegA<=FADDInstRegA[13:10];
	FADDDSTRegB<=FADDInstRegB[13:10];
	
	// FMUL channel
	FMULInstRegA<=FMULInstBusA;
	FMULInstRegB<=FMULInstBusB;
	FMULACTRegA<=FMULInstRegA[0];
	FMULACTRegB<=FMULInstRegB[0];

	FMULBypassARegA[0]<=FADDRDYRA & (FADDDSTRA==FMULInstBusA[4:1]);
	FMULBypassARegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FMULInstBusA[4:1]);
	FMULBypassARegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FMULInstBusA[4:1]);
	FMULBypassARegA[3]<=ALURDYRA & (ALUDSTRA==FMULInstBusA[4:1]);
	FMULBypassARegA[4]<=ShiftRDYR & (ShiftDSTR==FMULInstBusA[4:1]);
	FMULBypassARegA[5]<=MiscRDYR & (MiscDSTR==FMULInstBusA[4:1]);
	FMULBypassARegA[6]<=FADDRDYRB & (FADDDSTRB==FMULInstBusA[4:1]);
	FMULBypassARegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FMULInstBusA[4:1]);
	FMULBypassARegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FMULInstBusA[4:1]);
	FMULBypassARegA[9]<=ALURDYRB & (ALUDSTRB==FMULInstBusA[4:1]);

	FMULBypassARegB[0]<=FADDRDYRA & (FADDDSTRA==FMULInstBusB[4:1]);
	FMULBypassARegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FMULInstBusB[4:1]);
	FMULBypassARegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FMULInstBusB[4:1]);
	FMULBypassARegB[3]<=ALURDYRA & (ALUDSTRA==FMULInstBusB[4:1]);
	FMULBypassARegB[4]<=ShiftRDYR & (ShiftDSTR==FMULInstBusB[4:1]);
	FMULBypassARegB[5]<=MiscRDYR & (MiscDSTR==FMULInstBusB[4:1]);
	FMULBypassARegB[6]<=FADDRDYRB & (FADDDSTRB==FMULInstBusB[4:1]);
	FMULBypassARegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FMULInstBusB[4:1]);
	FMULBypassARegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FMULInstBusB[4:1]);
	FMULBypassARegB[9]<=ALURDYRB & (ALUDSTRB==FMULInstBusB[4:1]);

	FMULARegA<=(GPR[FMULInstRegA[4:1]] & {128{~(|FMULBypassARegA)}})|
				(FADDRA & {128{FMULBypassARegA[0]}}) |
				({64'd0, FMULRA & {64{FMULBypassARegA[1]}}}) |
				(FMULRQA & {128{FMULBypassARegA[2]}}) |
				({GPR[FMULInstRegA[4:1]][127:64], ALURA} & {128{FMULBypassARegA[3]}}) |
				({GPR[FMULInstRegA[4:1]][127:64], ShiftR} & {128{FMULBypassARegA[4]}}) |
				(MiscR & {128{FMULBypassARegA[5]}})|
				(FADDRB & {128{FMULBypassARegA[6]}}) |
				({64'd0, FMULRB & {64{FMULBypassARegA[7]}}}) |
				(FMULRQB & {128{FMULBypassARegA[8]}}) |
				({GPR[FMULInstRegA[4:1]][127:64], ALURB} & {128{FMULBypassARegA[9]}});

	FMULARegB<=(GPR[FMULInstRegB[4:1]] & {128{~(|FMULBypassARegB)}})|
				(FADDRA & {128{FMULBypassARegB[0]}}) |
				({64'd0, FMULRA & {64{FMULBypassARegB[1]}}}) |
				(FMULRQA & {128{FMULBypassARegB[2]}}) |
				({GPR[FMULInstRegB[4:1]][127:64], ALURA} & {128{FMULBypassARegB[3]}}) |
				({GPR[FMULInstRegB[4:1]][127:64], ShiftR} & {128{FMULBypassARegB[4]}}) |
				(MiscR & {128{FMULBypassARegB[5]}})|
				(FADDRB & {128{FMULBypassARegB[6]}}) |
				({64'd0, FMULRB & {64{FMULBypassARegB[7]}}}) |
				(FMULRQB & {128{FMULBypassARegB[8]}}) |
				({GPR[FMULInstRegB[4:1]][127:64], ALURB} & {128{FMULBypassARegB[9]}});

	FMULSARegA<=(AFR[FMULInstRegA[4:1]][24:22] & {3{~(|FMULBypassARegA)}})|
				(FADDSRA & {3{FMULBypassARegA[0]}})|
				({2'd1, FMULSRA} & {3{FMULBypassARegA[1]}})|
				({FMULBypassARegA[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FMULBypassARegA[3]}}})|
				({1'b0, ShiftSRReg & {2{FMULBypassARegA[4]}}})|
				(MiscSRReg & {3{FMULBypassARegA[5]}})|
				(FADDSRB & {3{FMULBypassARegA[6]}})|
				({2'd1, FMULSRB} & {3{FMULBypassARegA[7]}})|
				({FMULBypassARegA[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FMULBypassARegA[9]}}});

	FMULSARegB<=(AFR[FMULInstRegB[4:1]][24:22] & {3{~(|FMULBypassARegB)}})|
				(FADDSRA & {3{FMULBypassARegB[0]}})|
				({2'd1, FMULSRA} & {3{FMULBypassARegB[1]}})|
				({FMULBypassARegB[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FMULBypassARegB[3]}}})|
				({1'b0, ShiftSRReg & {2{FMULBypassARegB[4]}}})|
				(MiscSRReg & {3{FMULBypassARegB[5]}})|
				(FADDSRB & {3{FMULBypassARegB[6]}})|
				({2'd1, FMULSRB} & {3{FMULBypassARegB[7]}})|
				({FMULBypassARegB[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FMULBypassARegB[9]}}});

	FMULBypassBRegA[0]<=FADDRDYRA & (FADDDSTRA==FMULInstBusA[8:5]);
	FMULBypassBRegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FMULInstBusA[8:5]);
	FMULBypassBRegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FMULInstBusA[8:5]);
	FMULBypassBRegA[3]<=ALURDYRA & (ALUDSTRA==FMULInstBusA[8:5]);
	FMULBypassBRegA[4]<=ShiftRDYR & (ShiftDSTR==FMULInstBusA[8:5]);
	FMULBypassBRegA[5]<=MiscRDYR & (MiscDSTR==FMULInstBusA[8:5]);
	FMULBypassBRegA[6]<=FADDRDYRB & (FADDDSTRB==FMULInstBusA[8:5]);
	FMULBypassBRegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FMULInstBusA[8:5]);
	FMULBypassBRegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FMULInstBusA[8:5]);
	FMULBypassBRegA[9]<=ALURDYRB & (ALUDSTRB==FMULInstBusA[8:5]);

	FMULBypassBRegB[0]<=FADDRDYRA & (FADDDSTRA==FMULInstBusB[8:5]);
	FMULBypassBRegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FMULInstBusB[8:5]);
	FMULBypassBRegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FMULInstBusB[8:5]);
	FMULBypassBRegB[3]<=ALURDYRA & (ALUDSTRA==FMULInstBusB[8:5]);
	FMULBypassBRegB[4]<=ShiftRDYR & (ShiftDSTR==FMULInstBusB[8:5]);
	FMULBypassBRegB[5]<=MiscRDYR & (MiscDSTR==FMULInstBusB[8:5]);
	FMULBypassBRegB[6]<=FADDRDYRB & (FADDDSTRB==FMULInstBusB[8:5]);
	FMULBypassBRegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FMULInstBusB[8:5]);
	FMULBypassBRegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FMULInstBusB[8:5]);
	FMULBypassBRegB[9]<=ALURDYRB & (ALUDSTRB==FMULInstBusB[8:5]);

	FMULBRegA<=(GPR[FMULInstRegA[8:5]] & {128{~(|FMULBypassBRegA)}})|
				(FADDRA & {128{FMULBypassBRegA[0]}}) |
				({64'd0, FMULRA & {64{FMULBypassBRegA[1]}}}) |
				(FMULRQA & {128{FMULBypassBRegA[2]}}) |
				({GPR[FMULInstRegA[8:5]][127:64], ALURA} & {128{FMULBypassBRegA[3]}}) |
				({GPR[FMULInstRegA[8:5]][127:64], ShiftR} & {128{FMULBypassBRegA[4]}}) |
				(MiscR & {128{FMULBypassBRegA[5]}})|
				(FADDRB & {128{FMULBypassBRegA[6]}}) |
				({64'd0, FMULRB & {64{FMULBypassBRegA[7]}}}) |
				(FMULRQB & {128{FMULBypassBRegA[8]}}) |
				({GPR[FMULInstRegA[8:5]][127:64], ALURB} & {128{FMULBypassBRegA[9]}});

	FMULBRegB<=(GPR[FMULInstRegB[8:5]] & {128{~(|FMULBypassBRegB)}})|
				(FADDRA & {128{FMULBypassBRegB[0]}}) |
				({64'd0, FMULRA & {64{FMULBypassBRegB[1]}}}) |
				(FMULRQA & {128{FMULBypassBRegB[2]}}) |
				({GPR[FMULInstRegB[8:5]][127:64], ALURA} & {128{FMULBypassBRegB[3]}}) |
				({GPR[FMULInstRegB[8:5]][127:64], ShiftR} & {128{FMULBypassBRegB[4]}}) |
				(MiscR & {128{FMULBypassBRegB[5]}})|
				(FADDRB & {128{FMULBypassBRegB[6]}}) |
				({64'd0, FMULRB & {64{FMULBypassBRegB[7]}}}) |
				(FMULRQB & {128{FMULBypassBRegB[8]}}) |
				({GPR[FMULInstRegB[8:5]][127:64], ALURB} & {128{FMULBypassBRegB[9]}});

	FMULSBRegA<=(AFR[FMULInstRegA[8:5]][24:22] & {3{~(|FMULBypassBRegA)}})|
				(FADDSRA & {3{FMULBypassBRegA[0]}})|
				({2'd1, FMULSRA} & {3{FMULBypassBRegA[1]}})|
				({FMULBypassBRegA[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FMULBypassBRegA[3]}}})|
				({1'b0, ShiftSRReg & {2{FMULBypassBRegA[4]}}})|
				(MiscSRReg & {3{FMULBypassBRegA[5]}})|
				(FADDSRB & {3{FMULBypassBRegA[6]}})|
				({2'd1, FMULSRB} & {3{FMULBypassBRegA[7]}})|
				({FMULBypassBRegA[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FMULBypassBRegA[9]}}});

	FMULSBRegB<=(AFR[FMULInstRegB[8:5]][24:22] & {3{~(|FMULBypassBRegB)}})|
				(FADDSRA & {3{FMULBypassBRegB[0]}})|
				({2'd1, FMULSRA} & {3{FMULBypassBRegB[1]}})|
				({FMULBypassBRegB[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{FMULBypassBRegB[3]}}})|
				({1'b0, ShiftSRReg & {2{FMULBypassBRegB[4]}}})|
				(MiscSRReg & {3{FMULBypassBRegB[5]}})|
				(FADDSRB & {3{FMULBypassBRegB[6]}})|
				({2'd1, FMULSRB} & {3{FMULBypassBRegB[7]}})|
				({FMULBypassBRegB[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{FMULBypassBRegB[9]}}});

	FMULDSTRegA<=FMULInstRegA[12:9];
	FMULDSTRegB<=FMULInstRegB[12:9];

//=================================================================================================
//							FMULACC Channel
//0 - ACT, 3:1 - ctrlSel, 7:4 - DST, 11:8 - CtrlOffsetReg, 15:12 - DataOffsetReg, 18:16 - DataSel, 19 - CMD 0-FMULLACC/1-FFT
	FMULACCReg[0]<=(FMULACCReg[0] | FMULACCBus[0]) & (~FMULACCReg[0] | (FMULACCACTReg & ~FMULACCNEXT)) & RESET;
	if (~FMULACCReg[0]) FMULACCReg[19:1]<=FMULACCBus[19:1];
	
	FMULACCACTReg<=((FMULACCACTReg & ~FMULACCNEXT) | FMULACCReg[0]) & RESET;
	
	FFT32NEXTReg<=FFT32NEXT;
	
	FFTBypassReg[0]<=FADDRDYRA & (FADDDSTRA==FMULACCBus[7:4]);
	FFTBypassReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FMULACCBus[7:4]);
	FFTBypassReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FMULACCBus[7:4]);
	FFTBypassReg[3]<=ALURDYRA & (ALUDSTRA==FMULACCBus[7:4]);
	FFTBypassReg[4]<=ShiftRDYR & (ShiftDSTR==FMULACCBus[7:4]);
	FFTBypassReg[5]<=MiscRDYR & (MiscDSTR==FMULACCBus[7:4]);
	FFTBypassReg[6]<=FADDRDYRB & (FADDDSTRB==FMULACCBus[7:4]);
	FFTBypassReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FMULACCBus[7:4]);
	FFTBypassReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FMULACCBus[7:4]);
	FFTBypassReg[9]<=ALURDYRB & (ALUDSTRB==FMULACCBus[7:4]);

	FMULACCBypassControlOffsetReg[0]<=FADDRDYRA & (FADDDSTRA==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[3]<=ALURDYRA & (ALUDSTRA==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[4]<=ShiftRDYR & (ShiftDSTR==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[5]<=MiscRDYR & (MiscDSTR==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[6]<=FADDRDYRB & (FADDDSTRB==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FMULACCBus[11:8]);
	FMULACCBypassControlOffsetReg[9]<=ALURDYRB & (ALUDSTRB==FMULACCBus[11:8]);

	FMULACCBypassDataOffsetReg[0]<=FADDRDYRA & (FADDDSTRA==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[3]<=ALURDYRA & (ALUDSTRA==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[4]<=ShiftRDYR & (ShiftDSTR==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[5]<=MiscRDYR & (MiscDSTR==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[6]<=FADDRDYRB & (FADDDSTRB==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FMULACCBus[15:12]);
	FMULACCBypassDataOffsetReg[9]<=ALURDYRB & (ALUDSTRB==FMULACCBus[15:12]);

	if (FMULACCNEXT | ~FMULACCACTReg)
		begin
		FMULACCDSTReg<=FMULACCReg[7:4];
		FMULACCCtrlSelReg<=FMULACCReg[3:1];
		FMULACCDataSelReg<=FMULACCReg[18:16];
		
		FMULACCCMDReg<=FMULACCReg[19];
		
		FFTCtrlBaseReg<=ADR[{FMULACCReg[3:1],1'b0}][36:3];
		FFTDataBaseReg<=ADR[{FMULACCReg[18:16],1'b0}][36:3];
		FFTCtrlSelReg<=ADR[{FMULACCReg[3:1],1'b1}][31:0];
		FFTDataSelReg<=ADR[{FMULACCReg[18:16],1'b1}][31:0];
		
		FFTParReg<=(GPR[FMULACCReg[7:4]][4:0] & {5{~(|FFTBypassReg)}})|
					(FADDRA[4:0] & {5{FFTBypassReg[0]}}) |
					(FMULRA[4:0] & {5{FFTBypassReg[1]}}) |
					(FMULRQA[4:0] & {5{FFTBypassReg[2]}}) |
					(ALURA[4:0] & {5{FFTBypassReg[3]}}) |
					(ShiftR[4:0] & {5{FFTBypassReg[4]}}) |
					(MiscR[4:0] & {5{FFTBypassReg[5]}}) |
					(FADDRB[4:0] & {5{FFTBypassReg[6]}}) |
					(FMULRB[4:0] & {5{FFTBypassReg[7]}}) |
					(FMULRQB[4:0] & {5{FFTBypassReg[8]}}) |
					(ALURB[4:0] & {5{FFTBypassReg[9]}});
					
		FFTIndexReg<=(GPR[FMULACCReg[7:4]][50:32] & {19{~(|FFTBypassReg)}})|
					(FADDRA[50:32] & {19{FFTBypassReg[0]}}) |
					(FMULRA[50:32] & {19{FFTBypassReg[1]}}) |
					(FMULRQA[50:32] & {19{FFTBypassReg[2]}}) |
					(ALURA[50:32] & {19{FFTBypassReg[3]}}) |
					(ShiftR[50:32] & {19{FFTBypassReg[4]}}) |
					(MiscR[50:32] & {19{FFTBypassReg[5]}}) |
					(FADDRB[50:32] & {19{FFTBypassReg[6]}}) |
					(FMULRB[50:32] & {19{FFTBypassReg[7]}}) |
					(FMULRQB[50:32] & {19{FFTBypassReg[8]}}) |
					(ALURB[50:32] & {19{FFTBypassReg[9]}});
		
		FMULACCCtrlOffsetReg<=(GPR[FMULACCReg[11:8]][36:3] & {34{~(|FMULACCBypassControlOffsetReg)}})|
					(FADDRA[36:3] & {34{FMULACCBypassControlOffsetReg[0]}}) |
					(FMULRA[36:3] & {34{FMULACCBypassControlOffsetReg[1]}}) |
					(FMULRQA[36:3] & {34{FMULACCBypassControlOffsetReg[2]}}) |
					(ALURA[36:3] & {34{FMULACCBypassControlOffsetReg[3]}}) |
					(ShiftR[36:3] & {34{FMULACCBypassControlOffsetReg[4]}}) |
					(MiscR[36:3] & {34{FMULACCBypassControlOffsetReg[5]}})|
					(FADDRB[36:3] & {34{FMULACCBypassControlOffsetReg[6]}}) |
					(FMULRB[36:3] & {34{FMULACCBypassControlOffsetReg[7]}}) |
					(FMULRQB[36:3] & {34{FMULACCBypassControlOffsetReg[8]}}) |
					(ALURB[36:3] & {34{FMULACCBypassControlOffsetReg[9]}});
		
		FMULACCDataOffsetReg<=(GPR[FMULACCReg[15:12]][36:2] & {35{~(|FMULACCBypassDataOffsetReg)}})|
					(FADDRA[36:2] & {35{FMULACCBypassDataOffsetReg[0]}}) |
					(FMULRA[36:2] & {35{FMULACCBypassDataOffsetReg[1]}}) |
					(FMULRQA[36:2] & {35{FMULACCBypassDataOffsetReg[2]}}) |
					(ALURA[36:2] & {35{FMULACCBypassDataOffsetReg[3]}}) |
					(ShiftR[36:2] & {35{FMULACCBypassDataOffsetReg[4]}}) |
					(MiscR[36:2] & {35{FMULACCBypassDataOffsetReg[5]}})|
					(FADDRB[36:2] & {35{FMULACCBypassDataOffsetReg[6]}}) |
					(FMULRB[36:2] & {35{FMULACCBypassDataOffsetReg[7]}}) |
					(FMULRQB[36:2] & {35{FMULACCBypassDataOffsetReg[8]}}) |
					(ALURB[36:2] & {35{FMULACCBypassDataOffsetReg[9]}});
		end
	FMULACCDRDYFlag<=DRDY & (TAGi[7:1]==7'b1100000);

//=================================================================================================
//							FDIV channel
	
	
	FDIVInstReg[0]<=(FDIVInstReg[0] | FDIVInstBus[0]) & (~FDIVInstReg[0] | (FDIVACTReg & ~FDIVNEXT));
	if (~FDIVInstReg[0]) FDIVInstReg[13:1]<=FDIVInstBus[13:1];
	
	FDIVACTReg<=(FDIVACTReg & ~FDIVNEXT) | FDIVInstReg[0];

	FDIVBypassAReg[0]<=FADDRDYRA & (FADDDSTRA==FDIVInstBus[4:1]);
	FDIVBypassAReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FDIVInstBus[4:1]);
	FDIVBypassAReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FDIVInstBus[4:1]);
	FDIVBypassAReg[3]<=ALURDYRA & (ALUDSTRA==FDIVInstBus[4:1]);
	FDIVBypassAReg[4]<=ShiftRDYR & (ShiftDSTR==FDIVInstBus[4:1]);
	FDIVBypassAReg[5]<=MiscRDYR & (MiscDSTR==FDIVInstBus[4:1]);
	FDIVBypassAReg[6]<=FADDRDYRB & (FADDDSTRB==FDIVInstBus[4:1]);
	FDIVBypassAReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FDIVInstBus[4:1]);
	FDIVBypassAReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FDIVInstBus[4:1]);
	FDIVBypassAReg[9]<=ALURDYRB & (ALUDSTRB==FDIVInstBus[4:1]);

	FDIVBypassBReg[0]<=FADDRDYRA & (FADDDSTRA==FDIVInstBus[8:5]);
	FDIVBypassBReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==FDIVInstBus[8:5]);
	FDIVBypassBReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==FDIVInstBus[8:5]);
	FDIVBypassBReg[3]<=ALURDYRA & (ALUDSTRA==FDIVInstBus[8:5]);
	FDIVBypassBReg[4]<=ShiftRDYR & (ShiftDSTR==FDIVInstBus[8:5]);
	FDIVBypassBReg[5]<=MiscRDYR & (MiscDSTR==FDIVInstBus[8:5]);
	FDIVBypassBReg[6]<=FADDRDYRB & (FADDDSTRB==FDIVInstBus[8:5]);
	FDIVBypassBReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==FDIVInstBus[8:5]);
	FDIVBypassBReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==FDIVInstBus[8:5]);
	FDIVBypassBReg[9]<=ALURDYRB & (ALUDSTRB==FDIVInstBus[8:5]);

	if (FDIVNEXT | ~FDIVACTReg)
		begin
		FDIVAReg<=(GPR[FDIVInstReg[4:1]] & {128{~(|FDIVBypassAReg)}})|
					(FADDRA & {128{FDIVBypassAReg[0]}}) |
					({64'd0, FMULRA & {64{FDIVBypassAReg[1]}}}) |
					(FMULRQA & {128{FDIVBypassAReg[2]}}) |
					({GPR[FDIVInstReg[4:1]][127:64], ALURA} & {128{FDIVBypassAReg[3]}}) |
					({GPR[FDIVInstReg[4:1]][127:64], ShiftR} & {128{FDIVBypassAReg[4]}}) |
					(MiscR & {128{FDIVBypassAReg[5]}})|
					(FADDRB & {128{FDIVBypassAReg[6]}}) |
					({64'd0, FMULRB & {64{FDIVBypassAReg[7]}}}) |
					(FMULRQB & {128{FDIVBypassAReg[8]}}) |
					({GPR[FDIVInstReg[4:1]][127:64], ALURB} & {128{FDIVBypassAReg[9]}});

		FDIVSAReg<=(AFR[FDIVInstReg[4:1]][24:22] & {3{~(|FDIVBypassAReg)}})|
					(FADDSRA & {3{FDIVBypassAReg[0]}})|
					({2'd1, FMULSRA} & {3{FDIVBypassAReg[1]}})|
					({FDIVBypassAReg[2], 2'd0}) |
					({1'b0, ALUSRRegA & {2{FDIVBypassAReg[3]}}})|
					({1'b0, ShiftSRReg & {2{FDIVBypassAReg[4]}}})|
					(MiscSRReg & {3{FDIVBypassAReg[5]}})|
					(FADDSRB & {3{FDIVBypassAReg[6]}})|
					({2'd1, FMULSRB} & {3{FDIVBypassAReg[7]}})|
					({FDIVBypassAReg[8], 2'd0}) |
					({1'b0, ALUSRRegB & {2{FDIVBypassAReg[9]}}});

		FDIVBReg<=(GPR[FDIVInstReg[8:5]] & {128{~(|FDIVBypassBReg)}})|
					(FADDRA & {128{FDIVBypassBReg[0]}}) |
					({64'd0, FMULRA & {64{FDIVBypassBReg[1]}}}) |
					(FMULRQA & {128{FDIVBypassBReg[2]}}) |
					({GPR[FDIVInstReg[8:5]][127:64], ALURA} & {128{FDIVBypassBReg[3]}}) |
					({GPR[FDIVInstReg[8:5]][127:64], ShiftR} & {128{FDIVBypassBReg[4]}}) |
					(MiscR & {128{FDIVBypassBReg[5]}}) |
					(FADDRB & {128{FDIVBypassBReg[6]}}) |
					({64'd0, FMULRB & {64{FDIVBypassBReg[7]}}}) |
					(FMULRQB & {128{FDIVBypassBReg[8]}}) |
					({GPR[FDIVInstReg[8:5]][127:64], ALURB} & {128{FDIVBypassBReg[9]}});

		FDIVSBReg<=(AFR[FDIVInstReg[8:5]][24:22] & {3{~(|FDIVBypassBReg)}})|
					(FADDSRA & {3{FDIVBypassBReg[0]}})|
					({2'd1, FMULSRA} & {3{FDIVBypassBReg[1]}})|
					({FDIVBypassBReg[2], 2'd0}) |
					({1'b0, ALUSRRegA & {2{FDIVBypassBReg[3]}}})|
					({1'b0, ShiftSRReg & {2{FDIVBypassBReg[4]}}})|
					(MiscSRReg & {3{FDIVBypassBReg[5]}})|
					(FADDSRB & {3{FDIVBypassBReg[6]}})|
					({2'd1, FMULSRB} & {3{FDIVBypassBReg[7]}})|
					({FDIVBypassBReg[8], 2'd0}) |
					({1'b0, ALUSRRegB & {2{FDIVBypassBReg[9]}}});

		FDIVDSTReg<=FDIVInstReg[12:9];
		FDIVCMDReg<=FDIVInstReg[13];
		end

//=================================================================================================
// 							ALU channel

	ALUInstRegA<=ALUInstBusA;
	ALUInstRegB<=ALUInstBusB;
	ALUACTRegA<=ALUInstRegA[0];
	ALUACTRegB<=ALUInstRegB[0];
	ALUOpCODERegA<={ALUInstRegA[24], ALUInstRegA[2:1]};
	ALUOpCODERegB<={ALUInstRegB[24], ALUInstRegB[2:1]};

	ALUBypassARegA[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusA[6:3]);
	ALUBypassARegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusA[6:3]);
	ALUBypassARegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusA[6:3]);
	ALUBypassARegA[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusA[6:3]);
	ALUBypassARegA[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusA[6:3]);
	ALUBypassARegA[5]<=MiscRDYR & (MiscDSTR==ALUInstBusA[6:3]);
	ALUBypassARegA[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusA[6:3]);
	ALUBypassARegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusA[6:3]);
	ALUBypassARegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusA[6:3]);
	ALUBypassARegA[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusA[6:3]);

	ALUBypassARegB[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusB[6:3]);
	ALUBypassARegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusB[6:3]);
	ALUBypassARegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusB[6:3]);
	ALUBypassARegB[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusB[6:3]);
	ALUBypassARegB[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusB[6:3]);
	ALUBypassARegB[5]<=MiscRDYR & (MiscDSTR==ALUInstBusB[6:3]);
	ALUBypassARegB[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusB[6:3]);
	ALUBypassARegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusB[6:3]);
	ALUBypassARegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusB[6:3]);
	ALUBypassARegB[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusB[6:3]);

	ALUARegA<=ALUInstRegA[15] ? {58'd0, ALUInstRegA[8:3]} :
				((GPR[ALUInstRegA[6:3]][63:0] & {64{~(|ALUBypassARegA)}}) |
				(FADDRA[63:0] & {64{ALUBypassARegA[0]}}) |
				(FMULRA & {64{ALUBypassARegA[1]}}) |
				(FMULRQA[63:0] & {64{ALUBypassARegA[2]}}) |
				(ALURA & {64{ALUBypassARegA[3]}}) |
				(ShiftR & {64{ALUBypassARegA[4]}}) |
				(MiscR[63:0] & {64{ALUBypassARegA[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassARegA[6]}}) |
				(FMULRB & {64{ALUBypassARegA[7]}}) |
				(FMULRQB[63:0] & {64{ALUBypassARegA[8]}}) |
				(ALURB & {64{ALUBypassARegA[9]}}));

	ALUARegB<=ALUInstRegB[15] ? {58'd0, ALUInstRegB[8:3]} :
				((GPR[ALUInstRegB[6:3]][63:0] & {64{~(|ALUBypassARegB)}}) |
				(FADDRA[63:0] & {64{ALUBypassARegB[0]}}) |
				(FMULRA & {64{ALUBypassARegB[1]}}) |
				(FMULRQA[63:0] & {64{ALUBypassARegB[2]}}) |
				(ALURA & {64{ALUBypassARegB[3]}}) |
				(ShiftR & {64{ALUBypassARegB[4]}}) |
				(MiscR[63:0] & {64{ALUBypassARegB[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassARegB[6]}}) |
				(FMULRB & {64{ALUBypassARegB[7]}}) |
				(FMULRQB[63:0] & {64{ALUBypassARegB[8]}}) |
				(ALURB & {64{ALUBypassARegB[9]}}));

	ALUSARegA<=((AFR[ALUInstRegA[6:3]][23:22] & {2{~(|ALUBypassARegA)}}) |
					(FADDSRA[1:0] & {2{ALUBypassARegA[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassARegA[1]}}) |
					(ALUSRRegA & {2{ALUBypassARegA[3]}}) |
					(ShiftSRReg & {2{ALUBypassARegA[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassARegA[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassARegA[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassARegA[7]}}) |
					(ALUSRRegB & {2{ALUBypassARegA[9]}})) & {2{~ALUInstRegA[15]}};

	ALUSARegB<=((AFR[ALUInstRegB[6:3]][23:22] & {2{~(|ALUBypassARegB)}}) |
					(FADDSRA[1:0] & {2{ALUBypassARegB[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassARegB[1]}}) |
					(ALUSRRegA & {2{ALUBypassARegB[3]}}) |
					(ShiftSRReg & {2{ALUBypassARegB[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassARegB[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassARegB[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassARegB[7]}}) |
					(ALUSRRegB & {2{ALUBypassARegB[9]}})) & {2{~ALUInstRegB[15]}};

	ALUBypassBRegA[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusA[10:7]);
	ALUBypassBRegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusA[10:7]);
	ALUBypassBRegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusA[10:7]);
	ALUBypassBRegA[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusA[10:7]);
	ALUBypassBRegA[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusA[10:7]);
	ALUBypassBRegA[5]<=MiscRDYR & (MiscDSTR==ALUInstBusA[10:7]);
	ALUBypassBRegA[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusA[10:7]);
	ALUBypassBRegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusA[10:7]);
	ALUBypassBRegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusA[10:7]);
	ALUBypassBRegA[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusA[10:7]);

	ALUBypassBRegB[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusB[10:7]);
	ALUBypassBRegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusB[10:7]);
	ALUBypassBRegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusB[10:7]);
	ALUBypassBRegB[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusB[10:7]);
	ALUBypassBRegB[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusB[10:7]);
	ALUBypassBRegB[5]<=MiscRDYR & (MiscDSTR==ALUInstBusB[10:7]);
	ALUBypassBRegB[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusB[10:7]);
	ALUBypassBRegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusB[10:7]);
	ALUBypassBRegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusB[10:7]);
	ALUBypassBRegB[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusB[10:7]);

	ALUBRegA<=ALUInstRegA[15] ? {58'd0, ALUInstRegA[14:9]} :
				((GPR[ALUInstRegA[10:7]][63:0] & {64{~(|ALUBypassBRegA)}}) |
				(FADDRA[63:0] & {64{ALUBypassBRegA[0]}}) |
				(FMULRA & {64{ALUBypassBRegA[1]}}) | 
				(FMULRQA[63:0] & {64{ALUBypassBRegA[2]}}) |
				(ALURA & {64{ALUBypassBRegA[3]}}) |
				(ShiftR & {64{ALUBypassBRegA[4]}}) |
				(MiscR[63:0] & {64{ALUBypassBRegA[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassBRegA[6]}}) |
				(FMULRB & {64{ALUBypassBRegA[7]}}) | 
				(FMULRQB[63:0] & {64{ALUBypassBRegA[8]}}) |
				(ALURB & {64{ALUBypassBRegA[9]}}));

	ALUBRegB<=ALUInstRegB[15] ? {58'd0, ALUInstRegB[14:9]} :
				((GPR[ALUInstRegB[10:7]][63:0] & {64{~(|ALUBypassBRegB)}}) |
				(FADDRA[63:0] & {64{ALUBypassBRegB[0]}}) |
				(FMULRA & {64{ALUBypassBRegB[1]}}) | 
				(FMULRQA[63:0] & {64{ALUBypassBRegB[2]}}) |
				(ALURA & {64{ALUBypassBRegB[3]}}) |
				(ShiftR & {64{ALUBypassBRegB[4]}}) |
				(MiscR[63:0] & {64{ALUBypassBRegB[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassBRegB[6]}}) |
				(FMULRB & {64{ALUBypassBRegB[7]}}) | 
				(FMULRQB[63:0] & {64{ALUBypassBRegB[8]}}) |
				(ALURB & {64{ALUBypassBRegB[9]}}));

	ALUSBRegA<=((AFR[ALUInstRegA[10:7]][23:22] & {2{~(|ALUBypassBRegA)}}) |
					(FADDSRA[1:0] & {2{ALUBypassBRegA[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassBRegA[1]}}) | 
					(ALUSRRegA & {2{ALUBypassBRegA[3]}}) |
					(ShiftSRReg & {2{ALUBypassBRegA[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassBRegA[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassBRegA[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassBRegA[7]}}) | 
					(ALUSRRegB & {2{ALUBypassBRegA[9]}})) & {2{~ALUInstRegA[15]}};

	ALUSBRegB<=((AFR[ALUInstRegB[10:7]][23:22] & {2{~(|ALUBypassBRegB)}}) |
					(FADDSRA[1:0] & {2{ALUBypassBRegB[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassBRegB[1]}}) | 
					(ALUSRRegA & {2{ALUBypassBRegB[3]}}) |
					(ShiftSRReg & {2{ALUBypassBRegB[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassBRegB[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassBRegB[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassBRegB[7]}}) | 
					(ALUSRRegB & {2{ALUBypassBRegB[9]}})) & {2{~ALUInstRegB[15]}};

	ALUBypassCRegA[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusA[19:16]);
	ALUBypassCRegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusA[19:16]);
	ALUBypassCRegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusA[19:16]);
	ALUBypassCRegA[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusA[19:16]);
	ALUBypassCRegA[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusA[19:16]);
	ALUBypassCRegA[5]<=MiscRDYR & (MiscDSTR==ALUInstBusA[19:16]);
	ALUBypassCRegA[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusA[19:16]);
	ALUBypassCRegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusA[19:16]);
	ALUBypassCRegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusA[19:16]);
	ALUBypassCRegA[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusA[19:16]);

	ALUBypassCRegB[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusB[19:16]);
	ALUBypassCRegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusB[19:16]);
	ALUBypassCRegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusB[19:16]);
	ALUBypassCRegB[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusB[19:16]);
	ALUBypassCRegB[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusB[19:16]);
	ALUBypassCRegB[5]<=MiscRDYR & (MiscDSTR==ALUInstBusB[19:16]);
	ALUBypassCRegB[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusB[19:16]);
	ALUBypassCRegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusB[19:16]);
	ALUBypassCRegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusB[19:16]);
	ALUBypassCRegB[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusB[19:16]);

	ALUCRegA<=(GPR[ALUInstRegA[19:16]][63:0] & {64{~(|ALUBypassCRegA)}}) |
				(FADDRA[63:0] & {64{ALUBypassCRegA[0]}}) |
				(FMULRA & {64{ALUBypassCRegA[1]}}) |
				(FMULRQA[63:0] & {64{ALUBypassCRegA[2]}}) |
				(ALURA & {64{ALUBypassCRegA[3]}}) |
				(ShiftR & {64{ALUBypassCRegA[4]}}) |
				(MiscR[63:0] & {64{ALUBypassCRegA[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassCRegA[6]}}) |
				(FMULRB & {64{ALUBypassCRegA[7]}}) |
				(FMULRQB[63:0] & {64{ALUBypassCRegA[8]}}) |
				(ALURB & {64{ALUBypassCRegA[9]}});

	ALUCRegB<=(GPR[ALUInstRegB[19:16]][63:0] & {64{~(|ALUBypassCRegB)}}) |
				(FADDRA[63:0] & {64{ALUBypassCRegB[0]}}) |
				(FMULRA & {64{ALUBypassCRegB[1]}}) |
				(FMULRQA[63:0] & {64{ALUBypassCRegB[2]}}) |
				(ALURA & {64{ALUBypassCRegB[3]}}) |
				(ShiftR & {64{ALUBypassCRegB[4]}}) |
				(MiscR[63:0] & {64{ALUBypassCRegB[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassCRegB[6]}}) |
				(FMULRB & {64{ALUBypassCRegB[7]}}) |
				(FMULRQB[63:0] & {64{ALUBypassCRegB[8]}}) |
				(ALURB & {64{ALUBypassCRegB[9]}});

	ALUSCRegA<=((AFR[ALUInstRegA[19:16]][23:22] & {2{~(|ALUBypassCRegA)}}) |
					(FADDSRA[1:0] & {2{ALUBypassCRegA[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassCRegA[1]}}) |
					(ALUSRRegA & {2{ALUBypassCRegA[3]}}) |
					(ShiftSRReg & {2{ALUBypassCRegA[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassCRegA[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassCRegA[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassCRegA[7]}}) |
					(ALUSRRegB & {2{ALUBypassCRegA[9]}})) & {2{ALUInstRegA[24]}};

	ALUSCRegB<=((AFR[ALUInstRegB[19:16]][23:22] & {2{~(|ALUBypassCRegB)}}) |
					(FADDSRA[1:0] & {2{ALUBypassCRegB[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassCRegB[1]}}) |
					(ALUSRRegA & {2{ALUBypassCRegB[3]}}) |
					(ShiftSRReg & {2{ALUBypassCRegB[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassCRegB[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassCRegB[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassCRegB[7]}}) |
					(ALUSRRegB & {2{ALUBypassCRegB[9]}})) & {2{ALUInstRegB[24]}};

	ALUBypassDRegA[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusA[23:20]);
	ALUBypassDRegA[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusA[23:20]);
	ALUBypassDRegA[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusA[23:20]);
	ALUBypassDRegA[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusA[23:20]);
	ALUBypassDRegA[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusA[23:20]);
	ALUBypassDRegA[5]<=MiscRDYR & (MiscDSTR==ALUInstBusA[23:20]);
	ALUBypassDRegA[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusA[23:20]);
	ALUBypassDRegA[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusA[23:20]);
	ALUBypassDRegA[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusA[23:20]);
	ALUBypassDRegA[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusA[23:20]);

	ALUBypassDRegB[0]<=FADDRDYRA & (FADDDSTRA==ALUInstBusB[23:20]);
	ALUBypassDRegB[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ALUInstBusB[23:20]);
	ALUBypassDRegB[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ALUInstBusB[23:20]);
	ALUBypassDRegB[3]<=ALURDYRA & (ALUDSTRA==ALUInstBusB[23:20]);
	ALUBypassDRegB[4]<=ShiftRDYR & (ShiftDSTR==ALUInstBusB[23:20]);
	ALUBypassDRegB[5]<=MiscRDYR & (MiscDSTR==ALUInstBusB[23:20]);
	ALUBypassDRegB[6]<=FADDRDYRB & (FADDDSTRB==ALUInstBusB[23:20]);
	ALUBypassDRegB[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ALUInstBusB[23:20]);
	ALUBypassDRegB[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ALUInstBusB[23:20]);
	ALUBypassDRegB[9]<=ALURDYRB & (ALUDSTRB==ALUInstBusB[23:20]);

	ALUDRegA<=(GPR[ALUInstRegA[23:20]][63:0] & {64{~(|ALUBypassDRegA)}}) |
				(FADDRA[63:0] & {64{ALUBypassDRegA[0]}}) |
				(FMULRA & {64{ALUBypassDRegA[1]}}) |
				(FMULRQA[63:0] & {64{ALUBypassDRegA[2]}}) |
				(ALURA & {64{ALUBypassDRegA[3]}}) |
				(ShiftR & {64{ALUBypassDRegA[4]}}) |
				(MiscR[63:0] & {64{ALUBypassDRegA[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassDRegA[6]}}) |
				(FMULRB & {64{ALUBypassDRegA[7]}}) |
				(FMULRQB[63:0] & {64{ALUBypassDRegA[8]}}) |
				(ALURB & {64{ALUBypassDRegA[9]}});

	ALUDRegB<=(GPR[ALUInstRegB[23:20]][63:0] & {64{~(|ALUBypassDRegB)}}) |
				(FADDRA[63:0] & {64{ALUBypassDRegB[0]}}) |
				(FMULRA & {64{ALUBypassDRegB[1]}}) |
				(FMULRQA[63:0] & {64{ALUBypassDRegB[2]}}) |
				(ALURA & {64{ALUBypassDRegB[3]}}) |
				(ShiftR & {64{ALUBypassDRegB[4]}}) |
				(MiscR[63:0] & {64{ALUBypassDRegB[5]}}) |
				(FADDRB[63:0] & {64{ALUBypassDRegB[6]}}) |
				(FMULRB & {64{ALUBypassDRegB[7]}}) |
				(FMULRQB[63:0] & {64{ALUBypassDRegB[8]}}) |
				(ALURB & {64{ALUBypassDRegB[9]}});

	ALUSDRegA<=((AFR[ALUInstRegA[23:20]][23:22] & {2{~(|ALUBypassDRegA)}}) |
					(FADDSRA[1:0] & {2{ALUBypassDRegA[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassDRegA[1]}}) |
					(ALUSRRegA & {2{ALUBypassDRegA[3]}}) |
					(ShiftSRReg & {2{ALUBypassDRegA[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassDRegA[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassDRegA[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassDRegA[7]}}) |
					(ALUSRRegB & {2{ALUBypassDRegA[9]}})) & {2{ALUInstRegA[24]}};

	ALUSDRegB<=((AFR[ALUInstRegB[23:20]][23:22] & {2{~(|ALUBypassDRegB)}}) |
					(FADDSRA[1:0] & {2{ALUBypassDRegB[0]}}) |
					({1'b1, FMULSRA} & {2{ALUBypassDRegB[1]}}) |
					(ALUSRRegA & {2{ALUBypassDRegB[3]}}) |
					(ShiftSRReg & {2{ALUBypassDRegB[4]}}) |
					(MiscSRReg[1:0] & {2{ALUBypassDRegB[5]}}) |
					(FADDSRB[1:0] & {2{ALUBypassDRegB[6]}}) |
					({1'b1, FMULSRB} & {2{ALUBypassDRegB[7]}}) |
					(ALUSRRegB & {2{ALUBypassDRegB[9]}})) & {2{ALUInstRegB[24]}};

	ALUDSTRegA<=ALUInstRegA[24] ? ALUInstRegA[23:20] : ALUInstRegA[14:11];
	ALUDSTRegB<=ALUInstRegB[24] ? ALUInstRegB[23:20] : ALUInstRegB[14:11];

//=================================================================================================
//							Shifter channel

	ShiftInstReg<=ShiftInstBus;
	ShiftACTReg<=ShiftInstReg[0];

	ShiftBypassAReg[0]<=FADDRDYRA & (FADDDSTRA==ShiftInstBus[12:9]);
	ShiftBypassAReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ShiftInstBus[12:9]);
	ShiftBypassAReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ShiftInstBus[12:9]);
	ShiftBypassAReg[3]<=ALURDYRA & (ALUDSTRA==ShiftInstBus[12:9]);
	ShiftBypassAReg[4]<=ShiftRDYR & (ShiftDSTR==ShiftInstBus[12:9]);
	ShiftBypassAReg[5]<=MiscRDYR & (MiscDSTR==ShiftInstBus[12:9]);
	ShiftBypassAReg[6]<=FADDRDYRB & (FADDDSTRB==ShiftInstBus[12:9]);
	ShiftBypassAReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ShiftInstBus[12:9]);
	ShiftBypassAReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ShiftInstBus[12:9]);
	ShiftBypassAReg[9]<=ALURDYRB & (ALUDSTRB==ShiftInstBus[12:9]);

	ShiftAReg<=(GPR[ShiftInstReg[12:9]][63:0] & {64{~(|ShiftBypassAReg)}}) | 
				(FADDRA[63:0] & {64{ShiftBypassAReg[0]}}) |
				(FMULRA & {64{ShiftBypassAReg[1]}}) | 
				(FMULRQA[63:0] & {64{ShiftBypassAReg[2]}}) |
				(ALURA & {64{ShiftBypassAReg[3]}}) |
				(ShiftR & {64{ShiftBypassAReg[4]}}) |
				(MiscR[63:0] & {64{ShiftBypassAReg[5]}}) |
				(FADDRB[63:0] & {64{ShiftBypassAReg[6]}}) |
				(FMULRB & {64{ShiftBypassAReg[7]}}) | 
				(FMULRQB[63:0] & {64{ShiftBypassAReg[8]}}) |
				(ALURB & {64{ShiftBypassAReg[9]}});

	ShiftSAReg<=(AFR[ShiftInstReg[12:9]][23:22] & {2{~(|ShiftBypassAReg)}}) |
				(FADDSRA[1:0] & {2{ShiftBypassAReg[0]}}) |
				({1'b1, FMULSRA} & {2{ShiftBypassAReg[1]}}) |
				(ALUSRRegA & {2{ShiftBypassAReg[3]}}) |
				(ShiftSRReg & {2{ShiftBypassAReg[4]}}) |
				(MiscSRReg[1:0] & {2{ShiftBypassAReg[5]}}) |
				(FADDSRB[1:0] & {2{ShiftBypassAReg[6]}}) |
				({1'b1, FMULSRB} & {2{ShiftBypassAReg[7]}}) |
				(ALUSRRegB & {2{ShiftBypassAReg[9]}});

	ShiftBypassBReg[0]<=FADDRDYRA & (FADDDSTRA==ShiftInstBus[8:5]);
	ShiftBypassBReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==ShiftInstBus[8:5]);
	ShiftBypassBReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==ShiftInstBus[8:5]);
	ShiftBypassBReg[3]<=ALURDYRA & (ALUDSTRA==ShiftInstBus[8:5]);
	ShiftBypassBReg[4]<=ShiftRDYR & (ShiftDSTR==ShiftInstBus[8:5]);
	ShiftBypassBReg[5]<=MiscRDYR & (MiscDSTR==ShiftInstBus[8:5]);
	ShiftBypassBReg[6]<=FADDRDYRB & (FADDDSTRB==ShiftInstBus[8:5]);
	ShiftBypassBReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==ShiftInstBus[8:5]);
	ShiftBypassBReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==ShiftInstBus[8:5]);
	ShiftBypassBReg[9]<=ALURDYRB & (ALUDSTRB==ShiftInstBus[8:5]);

	ShiftBReg<=ShiftInstReg[4] ? ((GPR[ShiftInstReg[8:5]][5:0] & {6{~(|ShiftBypassBReg)}}) | 
								(FADDRA[5:0] & {6{ShiftBypassBReg[0]}}) |
								(FMULRA[5:0] & {6{ShiftBypassBReg[1]}}) | 
								(FMULRQA[5:0] & {6{ShiftBypassBReg[2]}}) |
								(ALURA[5:0] & {6{ShiftBypassBReg[3]}}) |
								(ShiftR[5:0] & {6{ShiftBypassBReg[4]}}) |
								(MiscR[5:0] & {6{ShiftBypassBReg[5]}}) |
								(FADDRB[5:0] & {6{ShiftBypassBReg[6]}}) |
								(FMULRB[5:0] & {6{ShiftBypassBReg[7]}}) | 
								(FMULRQB[5:0] & {6{ShiftBypassBReg[8]}}) |
								(ALURB[5:0] & {6{ShiftBypassBReg[9]}})) : {2'b00, ShiftInstReg[8:5]};							

	ShiftDSTReg<=ShiftInstReg[12:9];
	ShiftOPRReg<=ShiftInstReg[3:1];

//=================================================================================================
//							miscellaneous operations channel

	MiscInstReg<=MiscInstBus;
	MiscACTReg<=MiscInstReg[0];

	MiscBypassAReg[0]<=FADDRDYRA & (FADDDSTRA==MiscInstBus[7:4]);
	MiscBypassAReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==MiscInstBus[7:4]);
	MiscBypassAReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==MiscInstBus[7:4]);
	MiscBypassAReg[3]<=ALURDYRA & (ALUDSTRA==MiscInstBus[7:4]);
	MiscBypassAReg[4]<=ShiftRDYR & (ShiftDSTR==MiscInstBus[7:4]);
	MiscBypassAReg[5]<=MiscRDYR & (MiscDSTR==MiscInstBus[7:4]);
	MiscBypassAReg[6]<=FADDRDYRB & (FADDDSTRB==MiscInstBus[7:4]);
	MiscBypassAReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==MiscInstBus[7:4]);
	MiscBypassAReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==MiscInstBus[7:4]);
	MiscBypassAReg[9]<=ALURDYRB & (ALUDSTRB==MiscInstBus[7:4]);

	MiscBypassBReg[0]<=FADDRDYRA & (FADDDSTRA==MiscInstBus[11:8]);
	MiscBypassBReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==MiscInstBus[11:8]);
	MiscBypassBReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==MiscInstBus[11:8]);
	MiscBypassBReg[3]<=ALURDYRA & (ALUDSTRA==MiscInstBus[11:8]);
	MiscBypassBReg[4]<=ShiftRDYR & (ShiftDSTR==MiscInstBus[11:8]);
	MiscBypassBReg[5]<=MiscRDYR & (MiscDSTR==MiscInstBus[11:8]);
	MiscBypassBReg[6]<=FADDRDYRB & (FADDDSTRB==MiscInstBus[11:8]);
	MiscBypassBReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==MiscInstBus[11:8]);
	MiscBypassBReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==MiscInstBus[11:8]);
	MiscBypassBReg[9]<=ALURDYRB & (ALUDSTRB==MiscInstBus[11:8]);
	
	MiscCINReg<=(AFR[MiscInstReg[11:8]][15:0] & {16{~MiscBypassBReg[3] & ~MiscBypassBReg[9]}}) |
				(ALUCOUTA & {16{MiscBypassBReg[3]}}) | (ALUCOUTB & {16{MiscBypassBReg[9]}});

	MiscAReg<=(MiscInstReg[3] & (~MiscInstReg[2] | ~MiscInstReg[1])) ? ((GPR[MiscInstReg[7:4]] & {128{~(|MiscBypassAReg)}}) | 
																		(FADDRA & {128{MiscBypassAReg[0]}}) |
																		({64'd0, FMULRA & {64{MiscBypassAReg[1]}}}) |
																		(FMULRQA & {128{MiscBypassAReg[2]}}) |
																		({GPR[MiscInstReg[7:4]][127:64], ALURA} & {128{MiscBypassAReg[3]}}) |
																		({GPR[MiscInstReg[7:4]][127:64], ShiftR} & {128{MiscBypassAReg[4]}}) |
																		(MiscR & {128{MiscBypassAReg[5]}}) |
																		(FADDRB & {128{MiscBypassAReg[6]}}) |
																		({64'd0, FMULRB & {64{MiscBypassAReg[7]}}}) |
																		(FMULRQB & {128{MiscBypassAReg[8]}}) |
																		({GPR[MiscInstReg[7:4]][127:64], ALURB} & {128{MiscBypassAReg[9]}})) :
																		((GPR[MiscInstReg[11:8]] & {128{~(|MiscBypassBReg)}}) | 
																		(FADDRA & {128{MiscBypassBReg[0]}}) |
																		({64'd0, FMULRA & {64{MiscBypassBReg[1]}}}) |
																		(FMULRQA & {128{MiscBypassBReg[2]}}) |
																		({GPR[MiscInstReg[11:8]][127:64], ALURA} & {128{MiscBypassBReg[3]}}) |
																		({GPR[MiscInstReg[11:8]][127:64], ShiftR} & {128{MiscBypassBReg[4]}}) |
																		(MiscR & {128{MiscBypassBReg[5]}}) |
																		(FADDRB & {128{MiscBypassBReg[6]}}) |
																		({64'd0, FMULRB & {64{MiscBypassBReg[7]}}}) |
																		(FMULRQB & {128{MiscBypassBReg[8]}}) |
																		({GPR[MiscInstReg[11:8]][127:64], ALURB} & {128{MiscBypassBReg[9]}}));

	MiscSAReg<=(MiscInstReg[3] & (~MiscInstReg[2] | ~MiscInstReg[1])) ? ((AFR[MiscInstReg[7:4]][24:22] & {3{~(|MiscBypassAReg)}})|
																		(FADDSRA & {3{MiscBypassAReg[0]}})|
																		({2'd1, FMULSRA} & {3{MiscBypassAReg[1]}})|
																		({MiscBypassAReg[2], 2'd0}) |
																		({1'b0, ALUSRRegA & {2{MiscBypassAReg[3]}}})|
																		({1'b0, ShiftSRReg & {2{MiscBypassAReg[4]}}})|
																		(MiscSRReg & {3{MiscBypassAReg[5]}})|
																		(FADDSRB & {3{MiscBypassAReg[6]}})|
																		({2'd1, FMULSRB} & {3{MiscBypassAReg[7]}})|
																		({MiscBypassAReg[8], 2'd0}) |
																		({1'b0, ALUSRRegB & {2{MiscBypassAReg[9]}}})) :
																		((AFR[MiscInstReg[11:8]][24:22] & {3{~(|MiscBypassBReg)}})|
																		(FADDSRA & {3{MiscBypassBReg[0]}})|
																		({2'd1, FMULSRA} & {3{MiscBypassBReg[1]}})|
																		({MiscBypassBReg[2], 2'd0}) |
																		({1'b0, ALUSRRegA & {2{MiscBypassBReg[3]}}})|
																		({1'b0, ShiftSRReg & {2{MiscBypassBReg[4]}}})|
																		(MiscSRReg & {3{MiscBypassBReg[5]}})|
																		(FADDSRB & {3{MiscBypassBReg[6]}})|
																		({2'd1, FMULSRB} & {3{MiscBypassBReg[7]}})|
																		({MiscBypassBReg[8], 2'd0}) |
																		({1'b0, ALUSRRegB & {2{MiscBypassBReg[9]}}}));

	MiscSDReg<=(AFR[MiscInstReg[11:8]][24:22] & {3{~(|MiscBypassBReg)}})|
				(FADDSRA & {3{MiscBypassBReg[0]}})|
				({2'd1, FMULSRA} & {3{MiscBypassBReg[1]}})|
				({MiscBypassBReg[2], 2'd0}) |
				({1'b0, ALUSRRegA & {2{MiscBypassBReg[3]}}})|
				({1'b0, ShiftSRReg & {2{MiscBypassBReg[4]}}})|
				(MiscSRReg & {3{MiscBypassBReg[5]}})|
				(FADDSRB & {3{MiscBypassBReg[6]}})|
				({2'd1, FMULSRB} & {3{MiscBypassBReg[7]}})|
				({MiscBypassBReg[8], 2'd0}) |
				({1'b0, ALUSRRegB & {2{MiscBypassBReg[9]}}});

	MiscDSTReg<=MiscInstReg[11:8];
	MiscOPRReg<=MiscInstReg[3:1];
	
//=================================================================================================
//							loop instruction channel

	LoopInstReg<=LoopInstBus;

	LoopBypassReg[0]<=FADDRDYRA & (FADDDSTRA==LoopInstBus[15:12]);
	LoopBypassReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==LoopInstBus[15:12]);
	LoopBypassReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==LoopInstBus[15:12]);
	LoopBypassReg[3]<=ALURDYRA & (ALUDSTRA==LoopInstBus[15:12]);
	LoopBypassReg[4]<=ShiftRDYR & (ShiftDSTR==LoopInstBus[15:12]);
	LoopBypassReg[5]<=MiscRDYR & (MiscDSTR==LoopInstBus[15:12]);
	LoopBypassReg[6]<=FADDRDYRB & (FADDDSTRB==LoopInstBus[15:12]);
	LoopBypassReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==LoopInstBus[15:12]);
	LoopBypassReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==LoopInstBus[15:12]);
	LoopBypassReg[9]<=ALURDYRB & (ALUDSTRB==LoopInstBus[15:12]);
	
//=================================================================================================
//							prefetcher channel
	PrefInstReg<=PrefInstBus;

	PrefBypassReg[0]<=FADDRDYRA & (FADDDSTRA==PrefInstBus[16:13]);
	PrefBypassReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==PrefInstBus[16:13]);
	PrefBypassReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==PrefInstBus[16:13]);
	PrefBypassReg[3]<=ALURDYRA & (ALUDSTRA==PrefInstBus[16:13]);
	PrefBypassReg[4]<=ShiftRDYR & (ShiftDSTR==PrefInstBus[16:13]);
	PrefBypassReg[5]<=MiscRDYR & (MiscDSTR==PrefInstBus[16:13]);
	PrefBypassReg[6]<=FADDRDYRB & (FADDDSTRB==PrefInstBus[16:13]);
	PrefBypassReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==PrefInstBus[16:13]);
	PrefBypassReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==PrefInstBus[16:13]);
	PrefBypassReg[9]<=ALURDYRB & (ALUDSTRB==PrefInstBus[16:13]);
	
	PrefCCBypassReg[0]<=FADDRDYRA & (FADDDSTRA==PrefInstBus[8:5]);
	PrefCCBypassReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==PrefInstBus[8:5]);
	PrefCCBypassReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==PrefInstBus[8:5]);
	PrefCCBypassReg[3]<=ALURDYRA & (ALUDSTRA==PrefInstBus[8:5]);
	PrefCCBypassReg[4]<=ShiftRDYR & (ShiftDSTR==PrefInstBus[8:5]);
	PrefCCBypassReg[5]<=MiscRDYR & (MiscDSTR==PrefInstBus[8:5]);
	PrefCCBypassReg[6]<=FADDRDYRB & (FADDDSTRB==PrefInstBus[8:5]);
	PrefCCBypassReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==PrefInstBus[8:5]);
	PrefCCBypassReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==PrefInstBus[8:5]);
	PrefCCBypassReg[9]<=ALURDYRB & (ALUDSTRB==PrefInstBus[8:5]);
	
	// register movement operation
	MovInstReg<=MovInstBus;

	CopyBypassReg[0]<=FADDRDYRA & (FADDDSTRA==MovInstBus[10:7]);
	CopyBypassReg[1]<=FMULRDYRA[0] & (FMULDSTRA[0]==MovInstBus[10:7]);
	CopyBypassReg[2]<=FMULRDYRA[1] & (FMULDSTRA[1]==MovInstBus[10:7]);
	CopyBypassReg[3]<=ALURDYRA & (ALUDSTRA==MovInstBus[10:7]);
	CopyBypassReg[4]<=ShiftRDYR & (ShiftDSTR==MovInstBus[10:7]);
	CopyBypassReg[5]<=MiscRDYR & (MiscDSTR==MovInstBus[10:7]);
	CopyBypassReg[6]<=FADDRDYRB & (FADDDSTRB==MovInstBus[10:7]);
	CopyBypassReg[7]<=FMULRDYRB[0] & (FMULDSTRB[0]==MovInstBus[10:7]);
	CopyBypassReg[8]<=FMULRDYRB[1] & (FMULDSTRB[1]==MovInstBus[10:7]);
	CopyBypassReg[9]<=ALURDYRB & (ALUDSTRB==MovInstBus[10:7]);

	if (&MovInstReg[2:0]) 	begin
							// load immediate data mode
							case (AFR[MovInstReg[14:11]][31:28])
								4'h0: MovReg<={{120{MovInstReg[10]}},MovInstReg[10:3]};
								4'h1: MovReg<={{112{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][7:0]};
								4'h2: MovReg<={{104{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][15:0]};
								4'h3: MovReg<={{96{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][23:0]};
								4'h4: MovReg<={{88{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][31:0]};
								4'h5: MovReg<={{80{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][39:0]};
								4'h6: MovReg<={{72{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][47:0]};
								4'h7: MovReg<={{64{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][55:0]};
								4'h8: MovReg<={{56{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][63:0]};
								4'h9: MovReg<={{48{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][71:0]};
								4'hA: MovReg<={{40{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][79:0]};
								4'hB: MovReg<={{32{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][87:0]};
								4'hC: MovReg<={{24{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][95:0]};
								4'hD: MovReg<={{16{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][103:0]};
								4'hE: MovReg<={{8{MovInstReg[10]}},MovInstReg[10:3],GPR[MovInstReg[14:11]][111:0]};
								4'hF: MovReg<={MovInstReg[10:3],GPR[MovInstReg[14:11]][119:0]};
								endcase
							// size
							MovSR[0]<=(~AFR[MovInstReg[14:11]][31] & AFR[MovInstReg[14:11]][30])|
										(~AFR[MovInstReg[14:11]][31] & ~AFR[MovInstReg[14:11]][30] & ~AFR[MovInstReg[14:11]][29] & AFR[MovInstReg[14:11]][28]);
							MovSR[1]<=(AFR[MovInstReg[14:11]][30] | AFR[MovInstReg[14:11]][29]) & ~AFR[MovInstReg[14:11]][31];
							MovSR[2]<=AFR[MovInstReg[14:11]][31];
							end
			else begin
				if (MovInstReg[2:0]==3'b001)	begin
												// COPY operations
												MovReg<=(GPR[MovInstReg[10:7]] & {128{~(|CopyBypassReg)}}) | 
														(FADDRA & {128{CopyBypassReg[0]}}) |
														({64'd0, FMULRA & {64{CopyBypassReg[1]}}}) |
														(FMULRQA & {128{CopyBypassReg[2]}}) |
														({GPR[MovInstReg[10:7]][127:64], ALURA} & {128{CopyBypassReg[3]}}) |
														({GPR[MovInstReg[10:7]][127:64], ShiftR} & {128{CopyBypassReg[4]}}) |
														(MiscR & {128{CopyBypassReg[5]}}) |
														(FADDRB & {128{CopyBypassReg[6]}}) |
														({64'd0, FMULRB & {64{CopyBypassReg[7]}}}) |
														(FMULRQB & {128{CopyBypassReg[8]}}) |
														({GPR[MovInstReg[10:7]][127:64], ALURB} & {128{CopyBypassReg[9]}});
												MovSR<=(AFR[MovInstReg[10:7]][24:22] & {3{~(|CopyBypassReg)}})|
														(FADDSRA & {3{CopyBypassReg[0]}})|
														({2'd1, FMULSRA} & {3{CopyBypassReg[1]}})|
														({CopyBypassReg[2], 2'd0}) |
														({1'b0, ALUSRRegA & {2{CopyBypassReg[3]}}})|
														({1'b0, ShiftSRReg & {2{CopyBypassReg[4]}}})|
														(MiscSRReg & {3{CopyBypassReg[5]}})|
														(FADDSRB & {3{CopyBypassReg[6]}})|
														({2'd1, FMULSRB} & {3{CopyBypassReg[7]}})|
														({CopyBypassReg[8], 2'd0}) |
														({1'b0, ALUSRRegB & {2{CopyBypassReg[9]}}});
												end
										else if (MovInstReg[2:0]==3'b011) 
												begin
												if (MovInstReg[7]) AFR[MovInstReg[14:11]][27:25]<=MovInstReg[10:8];  // AMODE
															else	AFR[MovInstReg[14:11]][24:22]<=MovInstReg[10:8]; // SIZE
												end
				end

	//
	// Memory operations and address register 
	//
	if (~MemDelayFlag & ~MemFifoFullFlag) MemInstReg<=MemInstBus;

	MemDelayFlag<=~MemDelayFlag & MemInstBus[0] & ((FADDRDYRA & (FADDDSTRA==MemInstBus[15:12])) | (FADDRDYRB & (FADDDSTRB==MemInstBus[15:12])) |
					(FMULRDYRA[0] & (FMULDSTRA[0]==MemInstBus[15:12])) | (FMULRDYRB[0] & (FMULDSTRB[0]==MemInstBus[15:12])) |
					(FMULRDYRA[1] & (FMULDSTRA[1]==MemInstBus[15:12])) | (FMULRDYRB[1] & (FMULDSTRB[1]==MemInstBus[15:12])) | 
					(ALURDYRA & (ALUDSTRA==MemInstBus[15:12])) | (ALURDYRB & (ALUDSTRB==MemInstBus[15:12])) |
					(ShiftRDYR & (ShiftDSTR==MemInstBus[15:12])) | (MiscRDYR & (MiscDSTR==MemInstBus[15:12])) | 
					(FADDRDYRA & (FADDDSTRA==MemInstBus[11:8])) | (FADDRDYRB & (FADDDSTRB==MemInstBus[11:8])) |
					(FMULRDYRA[0] & (FMULDSTRA[0]==MemInstBus[11:8])) | (FMULRDYRB[0] & (FMULDSTRB[0]==MemInstBus[11:8])) |
					(FMULRDYRA[1] & (FMULDSTRA[1]==MemInstBus[11:8])) | (FMULRDYRB[1] & (FMULDSTRB[1]==MemInstBus[11:8])) |
					(ALURDYRA & (ALUDSTRA==MemInstBus[11:8])) | (ALURDYRB & (ALUDSTRB==MemInstBus[11:8])) |
					(ShiftRDYR & (ShiftDSTR==MemInstBus[11:8])) | (MiscRDYR & (MiscDSTR==MemInstBus[11:8])));	

	// busy flag of memory command
	MemBusy<=(MemBusy & ~MemLoadOffset & (~MemLoadSel | (MemDST=={CheckSEL,CheckACT})) & ~MemReadAR & ~(MemNext & ~FMULACCMemACT)) | MemCNT[1] | MemCNT[0] | ~MemFifoEmpty;
	
	// Memory interface unit operation flags
	if ((~MemBusy | (MemNext & ~FMULACCMemACT) | MemLoadOffset | (MemLoadSel & (MemDST!={CheckSEL,CheckACT})) | MemReadAR) & ~MemCNT[1] & ~MemCNT[0])
		begin
		// Read AR
		MemReadAR<=~MemFifoEmpty & ~MemFifoBus[3] & MemFifoBus[2] & ~MemFifoBus[1] & MemFifoBus[0] & ~MemFifoBus[215] & ~MemFifoBus[216];
		// Load AR (offset)
		MemLoadOffset<=~MemFifoEmpty & ~MemFifoBus[3] & MemFifoBus[2] & MemFifoBus[1] & ~MemFifoBus[0] & ~MemFifoBus[11] & ~MemFifoBus[215] & ~MemFifoBus[216];
		// Load AR (selector)
		MemLoadSel<=~MemFifoEmpty & ~MemFifoBus[3] & MemFifoBus[2] & MemFifoBus[1] & ~MemFifoBus[0] & MemFifoBus[11] & ~MemFifoBus[215] & ~MemFifoBus[216];
		// Request flag to the ATU
		MemReq<=~MemFifoEmpty & (MemFifoBus[3] | (~MemFifoBus[2] & ~MemFifoBus[1] & ~MemFifoBus[0]) |
												(MemFifoBus[2] & MemFifoBus[1] & MemFifoBus[0])) & ~MemFifoBus[215] & ~MemFifoBus[216];
		// Read/Write flag
		MemOpr<=MemFifoBus[3];
		// PUsh/POP/LDST flags
		MemPUSH<=~MemFifoEmpty & ~MemFifoBus[3] & MemFifoBus[2] & MemFifoBus[1] & MemFifoBus[0] & ~MemFifoBus[215] & ~MemFifoBus[216];
		MemPOP<=~MemFifoEmpty & MemFifoBus[3] & MemFifoBus[2] & MemFifoBus[1] & MemFifoBus[0] & ~MemFifoBus[215] & ~MemFifoBus[216];
		MemLDST<=~MemFifoEmpty & ((MemFifoBus[3] & (~MemFifoBus[2] | ~MemFifoBus[1] | ~MemFifoBus[0])) |
									(~MemFifoBus[3] & ~MemFifoBus[2] & ~MemFifoBus[1] & ~MemFifoBus[0])) & ~MemFifoBus[215] & ~MemFifoBus[216];
		MemLDO<=~MemFifoEmpty & MemFifoBus[3] & MemFifoBus[2] & ~MemFifoBus[1] & ~MemFifoBus[0] & ~MemFifoBus[215] & ~MemFifoBus[216];
		MemADRPushPop<=~MemFifoEmpty & MemFifoBus[2] & MemFifoBus[1] & MemFifoBus[0] & MemFifoBus[10] & ~MemFifoBus[215] & ~MemFifoBus[216];
		
		PrefCallReg<=~MemFifoEmpty & MemFifoBus[215];
		PrefRetReg<=~MemFifoEmpty & MemFifoBus[216];
		// Size
		if (MemFifoBus[3:0]==4'b0000) MemSize<=MemFifoBus[207:205];
								else MemSize<=MemFifoBus[2:0];
		// SEL field register
		if (MemFifoBus[3:0]==4'b0110) MemSEL<=MemFifoBus[14:12];
								else MemSEL<=MemFifoBus[6:4];
		// DST field register
		MemDST<=MemFifoBus[14:11];
		// Offset from GPR
		MemGPROffset<=MemFifoBus[51:15];
		// Offset register
		MemOFF<=MemFifoBus[10:7];
		// address mode
		MemAMode<=MemFifoBus[54:52];
		// GPR flags
		MemAFR<=MemFifoBus[214:183];
		// GPR
		MemGPR<=MemFifoBus[182:55];
		// data to GPR
		ARData<=ADR[MemOFF];
		end
	// Count of the bus cycles
	if ((~MemBusy | (MemNext & ~FMULACCMemACT) | MemLoadOffset | (MemLoadSel & (MemDST!={CheckSEL,CheckACT})) | MemReadAR) & ~MemFifoEmpty & (MemCNT==2'd0) & ~MemFifoBus[215] & ~MemFifoBus[216])
					begin
					MemCNT[0]<=(MemFifoBus[3:0]==4'b1100) |
							((MemFifoBus[3:0]==4'b0000) & MemFifoBus[207]);
					MemCNT[1]<=~MemFifoBus[10] & (MemFifoBus[2:0]==3'b111);
					end
				else if (MemNext & (MemCNT!=2'b00) & ~FMULACCMemACT) MemCNT<=MemCNT-2'd1;

	// resetting the descriptor valid flags 
	for (i=0; i<8; i=i+1)
		if (MemLoadSel & (MemSEL==i) & (MemDST!={CheckSEL,CheckACT & ~CheckAR[3]})) DTR[i][155]<=DTR[i][155] & (MemGPROffset[31:0]==ADR[{MemSEL,1'b1}][31:0]);
			else if (MemLSelNode & (TAGiReg[3:1]==i)) DTR[i][155]<=DTR[i][155] & (DTi[31:0]==ADR[TAGiReg[3:0]][31:0]);
	
	// second cycle for 128-bit transfers
	if ((MemNext & ~FMULACCMemACT) | ~MemBusy) MemSecondCycle<=(MemCNT==2'b01);
	//
	// processing address registers
	//
	for (i=0; i<16; i=i+1)
		if (i[0])
				begin
				// for selector registers
				if ((i!=15) & (i!=13))
						begin
						if (MemASelNode[i])	ADR[i]<=DTi[36:0];
							else if (MemLoadSel & (MemDST==i) & ((MemDST!={CheckSEL,CheckACT & ~CheckAR[3]}) | MemNext)) ADR[i]<=MemGPROffset;
						end
					else begin
						// stack selector and code selector can't be loaded from GPR's
						if (MemASelNode[i]) ADR[i]<=DTi[36:0];
							else if (MemLoadSel & (MemDST==i) & ~CPL[1] & ~CPL[0]) ADR[i]<=MemGPROffset;
						end
				end
			else begin
				// for offset registers
				if (i==14)
						begin
						// stack offset can be loaded from memory or modified in PUSH/POP/CALL/RET operations
						if (MemASelNode[i]) ADR[i]<=DTi[36:0];
							else if (MemLoadOffset & (MemDST==i)) ADR[i]<=MemGPROffset;
								else if ((MemPUSH | PrefCallReg) & MemNext & ~FMULACCMemACT) ADR[i]<=ADR[i]-8;
									else if ((MemPOP | PrefRetReg) & MemNext & ~FMULACCMemACT) ADR[i]<=ADR[i]+8;
						end
					else begin
						// all other offset registers
						if (MemASelNode[i]) ADR[i]<=DTi[36:0];
							else if (MemLoadOffset & (MemDST==i)) ADR[i]<=MemGPROffset;
									else if (MemLDST & MemNext & ~FMULACCMemACT & (({1'b0,MemSEL}<<1)==i) & MemReq & ~MemCNT[1] & ~MemCNT[0])
										begin
										if (MemAMode==3'b001) ADR[i]<=ADR[i]+MemGPROffset;
											else if (MemAMode[2] & ~MemAMode[0]) ADR[i]<=ADR[i]+MemoryOSValue;
												else if (MemAMode[2] & MemAMode[0]) ADR[i]<=ADR[i]-MemoryOSValue;
										end
						end
				end
	//
	// Conversion logical address to physical with access verification
	//
	CheckACT<=(CheckACT  & ~MemNext) | MemReq | PrefACT | PrefCallReg | PrefRetReg | FMULACCMemACT;
	
	// check offset and access type stage
	if (MemNext)
		begin
		// prefetcher flag
		CheckPref<=PrefACT & ~MemReq & ~PrefCallReg & ~PrefRetReg & ~FMULACCMemACT;
		// selector index
		if (FMULACCMemACT) CheckSEL<=FMULACCMemSEL;
			else if (PrefCallReg | PrefRetReg) CheckSEL<=3'd7;
					else if (MemReq) CheckSEL<=MemSEL | {3{MemPUSH | MemPOP}};
							else CheckSEL<=3'd6;

		// Command
		if (PrefCallReg) CheckCMD<=FMULACCMemACT;
			else if (MemReq) CheckCMD<=MemOpr | FMULACCMemACT | MemPOP;
					else CheckCMD<=1'b1;

		// operand size
		if (FMULACCMemACT) CheckOS<={1'b1,FMULACCSIZE};
			else if (MemReq) CheckOS<=MemSize[1:0] | {2{MemSize[2]}};
					else CheckOS<=2'b11;
		// Forming OFFSET 
		if (FMULACCMemACT) CheckOffset<=ADR[{1'b0,FMULACCMemSEL}<<1]+{FMULACCMemOffset,2'd0};
			else if (~MemReq & ~PrefCallReg & ~PrefRetReg) CheckOffset<=PrefOffset;
				else if (MemPUSH | PrefCallReg) CheckOffset<=ADR[14]-36'd8;
					else if (MemPOP | PrefRetReg) CheckOffset<=ADR[14];
							else case (MemAMode)
								3'b000 : CheckOffset<=ADR[{1'b0,MemSEL}<<1]+{33'd0,MemSecondCycle,3'd0};
								3'b001 : CheckOffset<=ADR[{1'b0,MemSEL}<<1]+{33'd0,MemSecondCycle,3'd0};
								3'b010 : CheckOffset<=MemGPROffset+{33'd0,MemSecondCycle,3'd0};
								3'b011 : CheckOffset<=ADR[{1'b0,MemSEL}<<1]+MemGPROffset+{33'd0,MemSecondCycle,3'd0};
								3'b100 : CheckOffset<=ADR[{1'b0,MemSEL}<<1]+{33'd0,MemSecondCycle,3'd0};
								3'b101 : CheckOffset<=ADR[{1'b0,MemSEL}<<1]+{33'd0,MemSecondCycle,3'd0};
								3'b110 : CheckOffset<=ADR[{1'b0,MemSEL}<<1]+MemGPROffset+{33'd0,MemSecondCycle,3'd0};
								3'b111 : CheckOffset<=ADR[{1'b0,MemSEL}<<1]+MemGPROffset+{33'd0,MemSecondCycle,3'd0};
								endcase
		// Base address limits and access rights
		if (FMULACCMemACT)
				begin
				CheckBase<=DTR[FMULACCMemSEL][39:0];
				CheckLL<=DTR[FMULACCMemSEL][71:40];
				CheckUL<=DTR[FMULACCMemSEL][103:72];
				CheckLowerSel<=DTR[FMULACCMemSEL][127:104];
				CheckUpperSel<=DTR[FMULACCMemSEL][151:128];
				CheckAR<=DTR[FMULACCMemSEL][155:152];
				CheckNetwork<=(CPU!=ADR[1+({1'b0,FMULACCMemSEL}<<1)][31:24]) & (|ADR[1+({1'b0,FMULACCMemSEL}<<1)][31:24]);
				CheckSelector<=ADR[1+({1'b0,FMULACCMemSEL}<<1)][31:0];
				end
			else begin
				if (MemPOP | MemPUSH | PrefCallReg | PrefRetReg)			//NEW
						begin
						// stack access
						CheckBase<=DTR[7][39:0];
						CheckLL<=DTR[7][71:40];
						CheckUL<=DTR[7][103:72];
						CheckLowerSel<=DTR[7][127:104];
						CheckUpperSel<=DTR[7][151:128];
						CheckAR<=DTR[7][155:152];
						CheckNetwork<=(CPU!=ADR[15][31:24]) & (|ADR[15][31:24]);
						CheckSelector<=ADR[15][31:0];
						end
					else begin
						if (MemReq)
							begin
							// data transactions
							CheckBase<=DTR[MemSEL][39:0];
							CheckLL<=DTR[MemSEL][71:40];
							CheckUL<=DTR[MemSEL][103:72];
							CheckLowerSel<=DTR[MemSEL][127:104];
							CheckUpperSel<=DTR[MemSEL][151:128];
							CheckAR<=DTR[MemSEL][155:152];
							CheckNetwork<=(CPU!=ADR[1+({1'b0,MemSEL}<<1)][31:24]) & (|ADR[1+({1'b0,MemSEL}<<1)][31:24]);
							CheckSelector<=ADR[1+({1'b0,MemSEL}<<1)][31:0];
							end
							else begin
							// code fetch
							CheckBase<=DTR[6][39:0];
							CheckLL<=DTR[6][71:40];
							CheckUL<=DTR[6][103:72];
							CheckLowerSel<=DTR[6][127:104];
							CheckUpperSel<=DTR[6][151:128];
							CheckAR<=DTR[6][155:152];
							CheckNetwork<=(CPU!=ADR[13][31:24]) & (|ADR[13][31:24]);
							CheckSelector<=ADR[13][31:0];
							end
					end
				end
		// forming data to memory
		if (PrefCallReg) CheckData<=MemGPR[63:0];
			else if (MemPUSH & (MemCNT==2'b10)) CheckData<=MemAFR;
					else if (MemPUSH & (MemCNT==2'b01)) CheckData<=MemGPR[127:64];
							else if (MemPUSH & MemSecondCycle) CheckData<=MemGPR[63:0];
									else if (MemPUSH & (MemCNT==2'b00)) CheckData<=ADR[MemDST];
											else if (MemSecondCycle) CheckData<=MemGPR[127:64];
													else CheckData<=MemGPR[63:0];
		// tag
		if (FMULACCMemACT) CheckTag<={7'b1100000, FMULACCTAGo};
			else if ((PrefCallReg | PrefRetReg) | (~MemReq & ~PrefCallReg & ~PrefRetReg))
						begin
						CheckTag[6:4]<=3'b110;
						CheckTag[3]<=PrefCallReg | PrefRetReg;
						CheckTag[2:0]<=PrefTag;
						CheckTag[7]<=1'b0;
						end
					else begin
						CheckTag[3:0]<=MemDST;
						CheckTag[4]<=(MemSecondCycle & MemLDST) | (~MemLDST & (MemCNT==2'b01)) | MemADRPushPop;
						CheckTag[5]<=(MemPUSH & (MemCNT==2'b10))|(MemPOP & (MemCNT==2'b00))| MemADRPushPop;
						CheckTag[6]<=1'b0;
						CheckTag[7]<=MemLDO;
						end
		end
	// reloading descriptor when he loaded from table
	if (DTRLoadedFlag)
		begin
		CheckBase<=DTR[CheckSEL][39:0];
		CheckLL<=DTR[CheckSEL][71:40];
		CheckUL<=DTR[CheckSEL][103:72];
		CheckLowerSel<=DTR[CheckSEL][127:104];
		CheckUpperSel<=DTR[CheckSEL][151:128];
		CheckAR<=DTR[CheckSEL][155:152];
		end

	//
	// output stage
	//
	// local memory access activation
	ACT<=(ACT & ~NEXT) | (CheckNext & CheckACT & CheckAR[3] & ~CheckNetwork & ~CheckAR[2] & (CheckOffset[36:5]>=CheckLL) & (CheckOffset[36:5]<CheckUL) & (CheckCMD | CheckAR[1]) & 
									(~CheckCMD | CheckAR[0])) | (DLMachine==LBS) | (DLMachine==LLSS) | (DLMachine==LSLS) |
									((DLMachine==STS) & CheckTag[6] & CheckTag[5] & ~CheckTag[4] & ~CheckTag[3]);
	// stream access activation
	StreamACT<=(StreamACT & ~StreamNEXT) | (CheckACT & CheckAR[3] & ~CheckNetwork & CheckAR[2] & CheckNext);
	
	// network access activation
	NetACT<=(NetACT & ~NetNEXT) | (CheckNext & CheckACT & CheckNetwork);
	
	if ((~ACT | NEXT) & (~StreamACT | StreamNEXT) & (~NetACT | NetNEXT))
		begin
		// command
		CMD<=CheckCMD | DescriptorLoadState;
		// operand size
		OS<=CheckOS | {2{DescriptorLoadState}};
		// forming physical address
		ADDRESS[2:0]<=DescriptorLoadState ? 3'b000 : CheckOffset[2:0];
		ADDRESS[3]<=DescriptorLoadState ? (DLMachine==LLSS) : CheckOffset[3];
		ADDRESS[4]<=DescriptorLoadState ? (DLMachine==LSLS) : CheckOffset[4];
		ADDRESS[44:5]<=DescriptorLoadState ? DTBASE + {16'd0, DLSelector} : (CheckNetwork ? {8'd0,CheckOffset[36:5]} : CheckBase+{8'd0,(CheckOffset[36:5]-CheckLL)});
		// offset
		OFFSET<=CheckOffset[36:0];
		// selector (for network accesses)
		SELECTOR<=CheckSelector;
		// data to memory
		DTo<=CheckData;
		// tag	
		TAGo[0]<=DescriptorLoadState ? (DLMachine==LLSS) : CheckTag[0];
		TAGo[1]<=DescriptorLoadState ? (DLMachine==LSLS) : CheckTag[1];
		TAGo[4:2]<=DescriptorLoadState ? CheckSEL : CheckTag[4:2] | {((DLMachine==STS) & CheckTag[6] & CheckTag[5] & ~CheckTag[4] & ~CheckTag[3]), 2'b00};
		TAGo[5]<=DescriptorLoadState ? 1'b0 : CheckTag[5];
		TAGo[6]<=DescriptorLoadState ? 1'b1 : CheckTag[6];
		TAGo[7]<=DescriptorLoadState ? 1'b0 : CheckTag[7];
		end

	//
	// Loading DT registers
	//
	DescriptorLoadState<=(DLMachine==CSS)|(DLMachine==LBS)|(DLMachine==LLSS)|(DLMachine==LSLS);
	// state machine for descriptor loading
		case (DLMachine)
				// wait state
				WS:	if (LoadNewDSC | LoadLowerDSC | LoadUpperDSC) DLMachine<=CSS;
						else if (AccessError) DLMachine<=AERSS;
								else DLMachine<=WS;
				// checking selector value
				CSS: if (DLSelector==24'd0) DLMachine<=ZSS;
						else if (DLSelector>=DTLIMIT) DLMachine<=INVSS;
							else DLMachine<=LBS;
				// load base address and access rights
				LBS: if (~ACT | NEXT) DLMachine<=LLSS;
						else DLMachine<=LBS;
				// load link selectors and check descriptor type
				LLSS: if (~ACT | NEXT) DLMachine<=LSLS;
						else DLMachine<=LLSS;
				// load segment limits
				LSLS: if (~ACT | NEXT) DLMachine<=RWS;
						else DLMachine<=LSLS;
				// waiting for transaction retry condition
				RWS: if (~RetryTransactionFlag) DLMachine<=RWS;
						else if (~ValidDescriptor) DLMachine<=INVOBS;
								else DLMachine<=WS;
				// zero selector reporting
				ZSS: DLMachine<=STS;
				// invalid selector reporting
				INVSS: DLMachine<=STS;
				// invalid object reporting (CPL or type)
				INVOBS: DLMachine<=STS;
				// access error
				AERSS: DLMachine<=STS;
				// skip transaction after error reporting
				STS: if (CheckTag[6] & CheckTag[5] & ~CheckTag[4] & ~CheckTag[3] & ~CheckNext) DLMachine<=STS;
						else DLMachine<=WS;
				endcase
	// temporary selector register
	if (DLMachine==WS) for (i=0; i<24; i=i+1) DLSelector[i]<=(LoadNewDSC & CheckSelector[i])|
															(LoadLowerDSC & CheckLowerSel[i])|
															(LoadUpperDSC & CheckUpperSel[i]);
				
	// 0 - base and AR, 1 - link selectors, 2 - limits
	for (i=0; i<8; i=i+1)
				if (DTRWriteFlag[i])
					case (TAGiReg[1:0])
						2'b00 : begin
								DTR[i][39:0]<=DTi[39:0];
								DTR[i][153:152]<=DTi[61:60];
								DTR[i][154]<=DTi[56];
								DTR[i][155]<=DTi[57] & (CPL<=DTi[59:58]) & ((TASKID==DTi[55:40]) | (~(|TASKID)) | (~(|DTi[55:40])));
								end
						2'b01 : begin
								DTR[i][127:104]<=DTi[23:0];
								DTR[i][151:128]<=DTi[55:32];
								end
						2'b10 :	begin
								DTR[i][103:40]<=DTi;
								end
						2'b11 :	DTR[i]<=156'hB000000000000FFFFFFFF000000000000000000;
						endcase
	DTRLoadedFlag<=DTRWriteFlag[8] & (TAGiReg[1:0]==2'b10);
	// flag to enable check transaction again
	RetryTransactionFlag<=DTRLoadedFlag;

	// valid descriptor flag
	if (DTRWriteFlag[8] & (TAGiReg[1:0]==2'b00))
		begin
		ValidDescriptor<=DTi[57] & (CPL<=DTi[59:58]) & ((TASKID==DTi[55:40]) | (~(|TASKID)) | (~(|DTi[55:40])));
		InvalidType<=~DTi[57];
		InvalidCPL<=(CPL>DTi[59:58]);
		InvalidTaskID<=(TASKID!=DTi[55:40]) & (|TASKID) & (|DTi[55:40]);
		InvalidSelector<=CheckSelector[23:0];
		end
	
	// skip read operation (validate flags)
	SkipDataRead<=CheckACT & CheckCMD & (DLMachine==STS) & ~CheckTag[6] & ~CheckTag[5];
	if (DLMachine==STS) STAGReg<=CheckTag[3:0];

	end

endmodule
